// hps_sub_sys.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module hps_sub_sys (
		input  wire         acp_0_clock_clk,                           //                  acp_0_clock.clk
		input  wire         acp_0_reset_reset,                         //                  acp_0_reset.reset
		input  wire         acp_0_csr_clock_clk,                       //              acp_0_csr_clock.clk
		input  wire         acp_0_csr_reset_reset,                     //              acp_0_csr_reset.reset
		input  wire         acp_0_csr_address,                         //                    acp_0_csr.address
		input  wire         acp_0_csr_read,                            //                             .read
		input  wire         acp_0_csr_write,                           //                             .write
		input  wire [31:0]  acp_0_csr_writedata,                       //                             .writedata
		output wire [31:0]  acp_0_csr_readdata,                        //                             .readdata
		input  wire [36:0]  acp_0_s0_araddr,                           //                     acp_0_s0.araddr
		input  wire [1:0]   acp_0_s0_arburst,                          //                             .arburst
		input  wire [3:0]   acp_0_s0_arcache,                          //                             .arcache
		input  wire [3:0]   acp_0_s0_arid,                             //                             .arid
		input  wire [7:0]   acp_0_s0_arlen,                            //                             .arlen
		input  wire         acp_0_s0_arlock,                           //                             .arlock
		input  wire [2:0]   acp_0_s0_arprot,                           //                             .arprot
		output wire         acp_0_s0_arready,                          //                             .arready
		input  wire [2:0]   acp_0_s0_arsize,                           //                             .arsize
		input  wire         acp_0_s0_arvalid,                          //                             .arvalid
		input  wire [36:0]  acp_0_s0_awaddr,                           //                             .awaddr
		input  wire [1:0]   acp_0_s0_awburst,                          //                             .awburst
		input  wire [3:0]   acp_0_s0_awcache,                          //                             .awcache
		input  wire [3:0]   acp_0_s0_awid,                             //                             .awid
		input  wire [7:0]   acp_0_s0_awlen,                            //                             .awlen
		input  wire         acp_0_s0_awlock,                           //                             .awlock
		input  wire [2:0]   acp_0_s0_awprot,                           //                             .awprot
		output wire         acp_0_s0_awready,                          //                             .awready
		input  wire [2:0]   acp_0_s0_awsize,                           //                             .awsize
		input  wire         acp_0_s0_awvalid,                          //                             .awvalid
		output wire [3:0]   acp_0_s0_bid,                              //                             .bid
		input  wire         acp_0_s0_bready,                           //                             .bready
		output wire [1:0]   acp_0_s0_bresp,                            //                             .bresp
		output wire         acp_0_s0_bvalid,                           //                             .bvalid
		output wire [511:0] acp_0_s0_rdata,                            //                             .rdata
		output wire [3:0]   acp_0_s0_rid,                              //                             .rid
		output wire         acp_0_s0_rlast,                            //                             .rlast
		input  wire         acp_0_s0_rready,                           //                             .rready
		output wire [1:0]   acp_0_s0_rresp,                            //                             .rresp
		output wire         acp_0_s0_rvalid,                           //                             .rvalid
		input  wire [511:0] acp_0_s0_wdata,                            //                             .wdata
		input  wire         acp_0_s0_wlast,                            //                             .wlast
		output wire         acp_0_s0_wready,                           //                             .wready
		input  wire [63:0]  acp_0_s0_wstrb,                            //                             .wstrb
		input  wire         acp_0_s0_wvalid,                           //                             .wvalid
		input  wire [43:0]  agilex_hps_f2h_stm_hw_events_stm_hwevents, // agilex_hps_f2h_stm_hw_events.stm_hwevents
		input  wire         agilex_hps_h2f_cs_ntrst,                   //            agilex_hps_h2f_cs.ntrst
		input  wire         agilex_hps_h2f_cs_tck,                     //                             .tck
		input  wire         agilex_hps_h2f_cs_tdi,                     //                             .tdi
		output wire         agilex_hps_h2f_cs_tdo,                     //                             .tdo
		output wire         agilex_hps_h2f_cs_tdoen,                   //                             .tdoen
		input  wire         agilex_hps_h2f_cs_tms,                     //                             .tms
		output wire         agilex_hps_hps_io_EMAC1_TX_CLK,            //            agilex_hps_hps_io.EMAC1_TX_CLK
		output wire         agilex_hps_hps_io_EMAC1_TXD0,              //                             .EMAC1_TXD0
		output wire         agilex_hps_hps_io_EMAC1_TXD1,              //                             .EMAC1_TXD1
		output wire         agilex_hps_hps_io_EMAC1_TXD2,              //                             .EMAC1_TXD2
		output wire         agilex_hps_hps_io_EMAC1_TXD3,              //                             .EMAC1_TXD3
		input  wire         agilex_hps_hps_io_EMAC1_RX_CTL,            //                             .EMAC1_RX_CTL
		output wire         agilex_hps_hps_io_EMAC1_TX_CTL,            //                             .EMAC1_TX_CTL
		input  wire         agilex_hps_hps_io_EMAC1_RX_CLK,            //                             .EMAC1_RX_CLK
		input  wire         agilex_hps_hps_io_EMAC1_RXD0,              //                             .EMAC1_RXD0
		input  wire         agilex_hps_hps_io_EMAC1_RXD1,              //                             .EMAC1_RXD1
		input  wire         agilex_hps_hps_io_EMAC1_RXD2,              //                             .EMAC1_RXD2
		input  wire         agilex_hps_hps_io_EMAC1_RXD3,              //                             .EMAC1_RXD3
		inout  wire         agilex_hps_hps_io_EMAC1_MDIO,              //                             .EMAC1_MDIO
		output wire         agilex_hps_hps_io_EMAC1_MDC,               //                             .EMAC1_MDC
		inout  wire         agilex_hps_hps_io_SDMMC_CMD,               //                             .SDMMC_CMD
		inout  wire         agilex_hps_hps_io_SDMMC_D0,                //                             .SDMMC_D0
		inout  wire         agilex_hps_hps_io_SDMMC_D1,                //                             .SDMMC_D1
		inout  wire         agilex_hps_hps_io_SDMMC_D2,                //                             .SDMMC_D2
		inout  wire         agilex_hps_hps_io_SDMMC_D3,                //                             .SDMMC_D3
		inout  wire         agilex_hps_hps_io_SDMMC_D4,                //                             .SDMMC_D4
		inout  wire         agilex_hps_hps_io_SDMMC_D5,                //                             .SDMMC_D5
		inout  wire         agilex_hps_hps_io_SDMMC_D6,                //                             .SDMMC_D6
		inout  wire         agilex_hps_hps_io_SDMMC_D7,                //                             .SDMMC_D7
		output wire         agilex_hps_hps_io_SDMMC_CCLK,              //                             .SDMMC_CCLK
		output wire         agilex_hps_hps_io_SPIM0_CLK,               //                             .SPIM0_CLK
		output wire         agilex_hps_hps_io_SPIM0_MOSI,              //                             .SPIM0_MOSI
		input  wire         agilex_hps_hps_io_SPIM0_MISO,              //                             .SPIM0_MISO
		output wire         agilex_hps_hps_io_SPIM0_SS0_N,             //                             .SPIM0_SS0_N
		output wire         agilex_hps_hps_io_SPIM1_CLK,               //                             .SPIM1_CLK
		output wire         agilex_hps_hps_io_SPIM1_MOSI,              //                             .SPIM1_MOSI
		input  wire         agilex_hps_hps_io_SPIM1_MISO,              //                             .SPIM1_MISO
		output wire         agilex_hps_hps_io_SPIM1_SS0_N,             //                             .SPIM1_SS0_N
		output wire         agilex_hps_hps_io_SPIM1_SS1_N,             //                             .SPIM1_SS1_N
		input  wire         agilex_hps_hps_io_UART1_RX,                //                             .UART1_RX
		output wire         agilex_hps_hps_io_UART1_TX,                //                             .UART1_TX
		inout  wire         agilex_hps_hps_io_I2C1_SDA,                //                             .I2C1_SDA
		inout  wire         agilex_hps_hps_io_I2C1_SCL,                //                             .I2C1_SCL
		input  wire         agilex_hps_hps_io_hps_osc_clk,             //                             .hps_osc_clk
		inout  wire         agilex_hps_hps_io_gpio0_io11,              //                             .gpio0_io11
		inout  wire         agilex_hps_hps_io_gpio0_io12,              //                             .gpio0_io12
		inout  wire         agilex_hps_hps_io_gpio0_io13,              //                             .gpio0_io13
		inout  wire         agilex_hps_hps_io_gpio0_io14,              //                             .gpio0_io14
		inout  wire         agilex_hps_hps_io_gpio0_io15,              //                             .gpio0_io15
		inout  wire         agilex_hps_hps_io_gpio0_io16,              //                             .gpio0_io16
		inout  wire         agilex_hps_hps_io_gpio0_io17,              //                             .gpio0_io17
		inout  wire         agilex_hps_hps_io_gpio0_io18,              //                             .gpio0_io18
		inout  wire         agilex_hps_hps_io_gpio1_io16,              //                             .gpio1_io16
		inout  wire         agilex_hps_hps_io_gpio1_io17,              //                             .gpio1_io17
		output wire         agilex_hps_h2f_reset_reset,                //         agilex_hps_h2f_reset.reset
		input  wire         agilex_hps_h2f_axi_clock_clk,              //     agilex_hps_h2f_axi_clock.clk
		input  wire         agilex_hps_h2f_axi_reset_reset_n,          //     agilex_hps_h2f_axi_reset.reset_n
		output wire [3:0]   agilex_hps_h2f_axi_master_awid,            //    agilex_hps_h2f_axi_master.awid
		output wire [31:0]  agilex_hps_h2f_axi_master_awaddr,          //                             .awaddr
		output wire [7:0]   agilex_hps_h2f_axi_master_awlen,           //                             .awlen
		output wire [2:0]   agilex_hps_h2f_axi_master_awsize,          //                             .awsize
		output wire [1:0]   agilex_hps_h2f_axi_master_awburst,         //                             .awburst
		output wire         agilex_hps_h2f_axi_master_awlock,          //                             .awlock
		output wire [3:0]   agilex_hps_h2f_axi_master_awcache,         //                             .awcache
		output wire [2:0]   agilex_hps_h2f_axi_master_awprot,          //                             .awprot
		output wire         agilex_hps_h2f_axi_master_awvalid,         //                             .awvalid
		input  wire         agilex_hps_h2f_axi_master_awready,         //                             .awready
		output wire [127:0] agilex_hps_h2f_axi_master_wdata,           //                             .wdata
		output wire [15:0]  agilex_hps_h2f_axi_master_wstrb,           //                             .wstrb
		output wire         agilex_hps_h2f_axi_master_wlast,           //                             .wlast
		output wire         agilex_hps_h2f_axi_master_wvalid,          //                             .wvalid
		input  wire         agilex_hps_h2f_axi_master_wready,          //                             .wready
		input  wire [3:0]   agilex_hps_h2f_axi_master_bid,             //                             .bid
		input  wire [1:0]   agilex_hps_h2f_axi_master_bresp,           //                             .bresp
		input  wire         agilex_hps_h2f_axi_master_bvalid,          //                             .bvalid
		output wire         agilex_hps_h2f_axi_master_bready,          //                             .bready
		output wire [3:0]   agilex_hps_h2f_axi_master_arid,            //                             .arid
		output wire [31:0]  agilex_hps_h2f_axi_master_araddr,          //                             .araddr
		output wire [7:0]   agilex_hps_h2f_axi_master_arlen,           //                             .arlen
		output wire [2:0]   agilex_hps_h2f_axi_master_arsize,          //                             .arsize
		output wire [1:0]   agilex_hps_h2f_axi_master_arburst,         //                             .arburst
		output wire         agilex_hps_h2f_axi_master_arlock,          //                             .arlock
		output wire [3:0]   agilex_hps_h2f_axi_master_arcache,         //                             .arcache
		output wire [2:0]   agilex_hps_h2f_axi_master_arprot,          //                             .arprot
		output wire         agilex_hps_h2f_axi_master_arvalid,         //                             .arvalid
		input  wire         agilex_hps_h2f_axi_master_arready,         //                             .arready
		input  wire [3:0]   agilex_hps_h2f_axi_master_rid,             //                             .rid
		input  wire [127:0] agilex_hps_h2f_axi_master_rdata,           //                             .rdata
		input  wire [1:0]   agilex_hps_h2f_axi_master_rresp,           //                             .rresp
		input  wire         agilex_hps_h2f_axi_master_rlast,           //                             .rlast
		input  wire         agilex_hps_h2f_axi_master_rvalid,          //                             .rvalid
		output wire         agilex_hps_h2f_axi_master_rready,          //                             .rready
		input  wire         agilex_hps_h2f_lw_axi_clock_clk,           //  agilex_hps_h2f_lw_axi_clock.clk
		input  wire         agilex_hps_h2f_lw_axi_reset_reset_n,       //  agilex_hps_h2f_lw_axi_reset.reset_n
		output wire [3:0]   agilex_hps_h2f_lw_axi_master_awid,         // agilex_hps_h2f_lw_axi_master.awid
		output wire [20:0]  agilex_hps_h2f_lw_axi_master_awaddr,       //                             .awaddr
		output wire [7:0]   agilex_hps_h2f_lw_axi_master_awlen,        //                             .awlen
		output wire [2:0]   agilex_hps_h2f_lw_axi_master_awsize,       //                             .awsize
		output wire [1:0]   agilex_hps_h2f_lw_axi_master_awburst,      //                             .awburst
		output wire         agilex_hps_h2f_lw_axi_master_awlock,       //                             .awlock
		output wire [3:0]   agilex_hps_h2f_lw_axi_master_awcache,      //                             .awcache
		output wire [2:0]   agilex_hps_h2f_lw_axi_master_awprot,       //                             .awprot
		output wire         agilex_hps_h2f_lw_axi_master_awvalid,      //                             .awvalid
		input  wire         agilex_hps_h2f_lw_axi_master_awready,      //                             .awready
		output wire [31:0]  agilex_hps_h2f_lw_axi_master_wdata,        //                             .wdata
		output wire [3:0]   agilex_hps_h2f_lw_axi_master_wstrb,        //                             .wstrb
		output wire         agilex_hps_h2f_lw_axi_master_wlast,        //                             .wlast
		output wire         agilex_hps_h2f_lw_axi_master_wvalid,       //                             .wvalid
		input  wire         agilex_hps_h2f_lw_axi_master_wready,       //                             .wready
		input  wire [3:0]   agilex_hps_h2f_lw_axi_master_bid,          //                             .bid
		input  wire [1:0]   agilex_hps_h2f_lw_axi_master_bresp,        //                             .bresp
		input  wire         agilex_hps_h2f_lw_axi_master_bvalid,       //                             .bvalid
		output wire         agilex_hps_h2f_lw_axi_master_bready,       //                             .bready
		output wire [3:0]   agilex_hps_h2f_lw_axi_master_arid,         //                             .arid
		output wire [20:0]  agilex_hps_h2f_lw_axi_master_araddr,       //                             .araddr
		output wire [7:0]   agilex_hps_h2f_lw_axi_master_arlen,        //                             .arlen
		output wire [2:0]   agilex_hps_h2f_lw_axi_master_arsize,       //                             .arsize
		output wire [1:0]   agilex_hps_h2f_lw_axi_master_arburst,      //                             .arburst
		output wire         agilex_hps_h2f_lw_axi_master_arlock,       //                             .arlock
		output wire [3:0]   agilex_hps_h2f_lw_axi_master_arcache,      //                             .arcache
		output wire [2:0]   agilex_hps_h2f_lw_axi_master_arprot,       //                             .arprot
		output wire         agilex_hps_h2f_lw_axi_master_arvalid,      //                             .arvalid
		input  wire         agilex_hps_h2f_lw_axi_master_arready,      //                             .arready
		input  wire [3:0]   agilex_hps_h2f_lw_axi_master_rid,          //                             .rid
		input  wire [31:0]  agilex_hps_h2f_lw_axi_master_rdata,        //                             .rdata
		input  wire [1:0]   agilex_hps_h2f_lw_axi_master_rresp,        //                             .rresp
		input  wire         agilex_hps_h2f_lw_axi_master_rlast,        //                             .rlast
		input  wire         agilex_hps_h2f_lw_axi_master_rvalid,       //                             .rvalid
		output wire         agilex_hps_h2f_lw_axi_master_rready,       //                             .rready
		input  wire         agilex_hps_f2h_axi_clock_clk,              //     agilex_hps_f2h_axi_clock.clk
		input  wire         agilex_hps_f2h_axi_reset_reset_n,          //     agilex_hps_f2h_axi_reset.reset_n
		input  wire [31:0]  agilex_hps_f2h_irq0_irq,                   //          agilex_hps_f2h_irq0.irq
		input  wire [31:0]  agilex_hps_f2h_irq1_irq,                   //          agilex_hps_f2h_irq1.irq
		input  wire         emif_hps_pll_ref_clk_clk,                  //         emif_hps_pll_ref_clk.clk
		input  wire         emif_hps_oct_oct_rzqin,                    //                 emif_hps_oct.oct_rzqin
		output wire [0:0]   emif_hps_mem_mem_ck,                       //                 emif_hps_mem.mem_ck
		output wire [0:0]   emif_hps_mem_mem_ck_n,                     //                             .mem_ck_n
		output wire [16:0]  emif_hps_mem_mem_a,                        //                             .mem_a
		output wire [0:0]   emif_hps_mem_mem_act_n,                    //                             .mem_act_n
		output wire [1:0]   emif_hps_mem_mem_ba,                       //                             .mem_ba
		output wire [0:0]   emif_hps_mem_mem_bg,                       //                             .mem_bg
		output wire [0:0]   emif_hps_mem_mem_cke,                      //                             .mem_cke
		output wire [1:0]   emif_hps_mem_mem_cs_n,                     //                             .mem_cs_n
		output wire [0:0]   emif_hps_mem_mem_odt,                      //                             .mem_odt
		output wire [0:0]   emif_hps_mem_mem_reset_n,                  //                             .mem_reset_n
		output wire [0:0]   emif_hps_mem_mem_par,                      //                             .mem_par
		input  wire [0:0]   emif_hps_mem_mem_alert_n,                  //                             .mem_alert_n
		inout  wire [8:0]   emif_hps_mem_mem_dqs,                      //                             .mem_dqs
		inout  wire [8:0]   emif_hps_mem_mem_dqs_n,                    //                             .mem_dqs_n
		inout  wire [71:0]  emif_hps_mem_mem_dq,                       //                             .mem_dq
		inout  wire [8:0]   emif_hps_mem_mem_dbi_n                     //                             .mem_dbi_n
	);

	wire     [1:0] agilex_axi_bridge_for_acp_0_m0_awburst;     // agilex_axi_bridge_for_acp_0:axm_m0_awburst -> agilex_hps:f2h_AWBURST
	wire     [7:0] agilex_axi_bridge_for_acp_0_m0_arlen;       // agilex_axi_bridge_for_acp_0:axm_m0_arlen -> agilex_hps:f2h_ARLEN
	wire     [3:0] agilex_axi_bridge_for_acp_0_m0_arqos;       // agilex_axi_bridge_for_acp_0:axm_m0_arqos -> agilex_hps:f2h_ARQOS
	wire    [22:0] agilex_axi_bridge_for_acp_0_m0_awuser;      // agilex_axi_bridge_for_acp_0:axm_m0_awuser -> agilex_hps:f2h_AWUSER
	wire     [3:0] agilex_axi_bridge_for_acp_0_m0_arsnoop;     // agilex_axi_bridge_for_acp_0:axm_m0_arsnoop -> agilex_hps:f2h_ARSNOOP
	wire           agilex_axi_bridge_for_acp_0_m0_wready;      // agilex_hps:f2h_WREADY -> agilex_axi_bridge_for_acp_0:axm_m0_wready
	wire    [63:0] agilex_axi_bridge_for_acp_0_m0_wstrb;       // agilex_axi_bridge_for_acp_0:axm_m0_wstrb -> agilex_hps:f2h_WSTRB
	wire     [2:0] agilex_axi_bridge_for_acp_0_m0_awsnoop;     // agilex_axi_bridge_for_acp_0:axm_m0_awsnoop -> agilex_hps:f2h_AWSNOOP
	wire     [4:0] agilex_axi_bridge_for_acp_0_m0_rid;         // agilex_hps:f2h_RID -> agilex_axi_bridge_for_acp_0:axm_m0_rid
	wire     [1:0] agilex_axi_bridge_for_acp_0_m0_arbar;       // agilex_axi_bridge_for_acp_0:axm_m0_arbar -> agilex_hps:f2h_ARBAR
	wire           agilex_axi_bridge_for_acp_0_m0_rready;      // agilex_axi_bridge_for_acp_0:axm_m0_rready -> agilex_hps:f2h_RREADY
	wire     [7:0] agilex_axi_bridge_for_acp_0_m0_awlen;       // agilex_axi_bridge_for_acp_0:axm_m0_awlen -> agilex_hps:f2h_AWLEN
	wire     [3:0] agilex_axi_bridge_for_acp_0_m0_awqos;       // agilex_axi_bridge_for_acp_0:axm_m0_awqos -> agilex_hps:f2h_AWQOS
	wire     [1:0] agilex_axi_bridge_for_acp_0_m0_awbar;       // agilex_axi_bridge_for_acp_0:axm_m0_awbar -> agilex_hps:f2h_AWBAR
	wire     [3:0] agilex_axi_bridge_for_acp_0_m0_arcache;     // agilex_axi_bridge_for_acp_0:axm_m0_arcache -> agilex_hps:f2h_ARCACHE
	wire    [36:0] agilex_axi_bridge_for_acp_0_m0_araddr;      // agilex_axi_bridge_for_acp_0:axm_m0_araddr -> agilex_hps:f2h_ARADDR
	wire           agilex_axi_bridge_for_acp_0_m0_wvalid;      // agilex_axi_bridge_for_acp_0:axm_m0_wvalid -> agilex_hps:f2h_WVALID
	wire     [2:0] agilex_axi_bridge_for_acp_0_m0_arprot;      // agilex_axi_bridge_for_acp_0:axm_m0_arprot -> agilex_hps:f2h_ARPROT
	wire           agilex_axi_bridge_for_acp_0_m0_arvalid;     // agilex_axi_bridge_for_acp_0:axm_m0_arvalid -> agilex_hps:f2h_ARVALID
	wire     [2:0] agilex_axi_bridge_for_acp_0_m0_awprot;      // agilex_axi_bridge_for_acp_0:axm_m0_awprot -> agilex_hps:f2h_AWPROT
	wire   [511:0] agilex_axi_bridge_for_acp_0_m0_wdata;       // agilex_axi_bridge_for_acp_0:axm_m0_wdata -> agilex_hps:f2h_WDATA
	wire     [4:0] agilex_axi_bridge_for_acp_0_m0_arid;        // agilex_axi_bridge_for_acp_0:axm_m0_arid -> agilex_hps:f2h_ARID
	wire     [3:0] agilex_axi_bridge_for_acp_0_m0_awcache;     // agilex_axi_bridge_for_acp_0:axm_m0_awcache -> agilex_hps:f2h_AWCACHE
	wire           agilex_axi_bridge_for_acp_0_m0_arlock;      // agilex_axi_bridge_for_acp_0:axm_m0_arlock -> agilex_hps:f2h_ARLOCK
	wire           agilex_axi_bridge_for_acp_0_m0_awlock;      // agilex_axi_bridge_for_acp_0:axm_m0_awlock -> agilex_hps:f2h_AWLOCK
	wire    [36:0] agilex_axi_bridge_for_acp_0_m0_awaddr;      // agilex_axi_bridge_for_acp_0:axm_m0_awaddr -> agilex_hps:f2h_AWADDR
	wire           agilex_axi_bridge_for_acp_0_m0_arready;     // agilex_hps:f2h_ARREADY -> agilex_axi_bridge_for_acp_0:axm_m0_arready
	wire     [1:0] agilex_axi_bridge_for_acp_0_m0_bresp;       // agilex_hps:f2h_BRESP -> agilex_axi_bridge_for_acp_0:axm_m0_bresp
	wire   [511:0] agilex_axi_bridge_for_acp_0_m0_rdata;       // agilex_hps:f2h_RDATA -> agilex_axi_bridge_for_acp_0:axm_m0_rdata
	wire     [1:0] agilex_axi_bridge_for_acp_0_m0_arburst;     // agilex_axi_bridge_for_acp_0:axm_m0_arburst -> agilex_hps:f2h_ARBURST
	wire           agilex_axi_bridge_for_acp_0_m0_awready;     // agilex_hps:f2h_AWREADY -> agilex_axi_bridge_for_acp_0:axm_m0_awready
	wire     [2:0] agilex_axi_bridge_for_acp_0_m0_arsize;      // agilex_axi_bridge_for_acp_0:axm_m0_arsize -> agilex_hps:f2h_ARSIZE
	wire           agilex_axi_bridge_for_acp_0_m0_bready;      // agilex_axi_bridge_for_acp_0:axm_m0_bready -> agilex_hps:f2h_BREADY
	wire           agilex_axi_bridge_for_acp_0_m0_rlast;       // agilex_hps:f2h_RLAST -> agilex_axi_bridge_for_acp_0:axm_m0_rlast
	wire     [1:0] agilex_axi_bridge_for_acp_0_m0_awdomain;    // agilex_axi_bridge_for_acp_0:axm_m0_awdomain -> agilex_hps:f2h_AWDOMAIN
	wire           agilex_axi_bridge_for_acp_0_m0_wlast;       // agilex_axi_bridge_for_acp_0:axm_m0_wlast -> agilex_hps:f2h_WLAST
	wire     [1:0] agilex_axi_bridge_for_acp_0_m0_ardomain;    // agilex_axi_bridge_for_acp_0:axm_m0_ardomain -> agilex_hps:f2h_ARDOMAIN
	wire     [1:0] agilex_axi_bridge_for_acp_0_m0_rresp;       // agilex_hps:f2h_RRESP -> agilex_axi_bridge_for_acp_0:axm_m0_rresp
	wire     [4:0] agilex_axi_bridge_for_acp_0_m0_awid;        // agilex_axi_bridge_for_acp_0:axm_m0_awid -> agilex_hps:f2h_AWID
	wire     [4:0] agilex_axi_bridge_for_acp_0_m0_bid;         // agilex_hps:f2h_BID -> agilex_axi_bridge_for_acp_0:axm_m0_bid
	wire           agilex_axi_bridge_for_acp_0_m0_bvalid;      // agilex_hps:f2h_BVALID -> agilex_axi_bridge_for_acp_0:axm_m0_bvalid
	wire    [22:0] agilex_axi_bridge_for_acp_0_m0_aruser;      // agilex_axi_bridge_for_acp_0:axm_m0_aruser -> agilex_hps:f2h_ARUSER
	wire     [2:0] agilex_axi_bridge_for_acp_0_m0_awsize;      // agilex_axi_bridge_for_acp_0:axm_m0_awsize -> agilex_hps:f2h_AWSIZE
	wire           agilex_axi_bridge_for_acp_0_m0_awvalid;     // agilex_axi_bridge_for_acp_0:axm_m0_awvalid -> agilex_hps:f2h_AWVALID
	wire           agilex_axi_bridge_for_acp_0_m0_rvalid;      // agilex_hps:f2h_RVALID -> agilex_axi_bridge_for_acp_0:axm_m0_rvalid
	wire           emif_calbus_0_emif_calbus_clk_clk;          // emif_calbus_0:calbus_clk -> emif_hps:calbus_clk
	wire    [31:0] emif_calbus_0_emif_calbus_0_calbus_wdata;   // emif_calbus_0:calbus_wdata_0 -> emif_hps:calbus_wdata
	wire    [19:0] emif_calbus_0_emif_calbus_0_calbus_address; // emif_calbus_0:calbus_address_0 -> emif_hps:calbus_address
	wire  [4095:0] emif_hps_emif_calbus_calbus_seq_param_tbl;  // emif_hps:calbus_seq_param_tbl -> emif_calbus_0:calbus_seq_param_tbl_0
	wire           emif_calbus_0_emif_calbus_0_calbus_read;    // emif_calbus_0:calbus_read_0 -> emif_hps:calbus_read
	wire           emif_calbus_0_emif_calbus_0_calbus_write;   // emif_calbus_0:calbus_write_0 -> emif_hps:calbus_write
	wire    [31:0] emif_hps_emif_calbus_calbus_rdata;          // emif_hps:calbus_rdata -> emif_calbus_0:calbus_rdata_0
	wire     [1:0] agilex_hps_hps_emif_gp_to_emif;             // agilex_hps:hps_emif_gp_to_emif -> emif_hps:hps_to_emif_gp
	wire  [4095:0] emif_hps_hps_emif_emif_to_hps;              // emif_hps:emif_to_hps -> agilex_hps:hps_emif_emif_to_hps
	wire     [0:0] emif_hps_hps_emif_emif_to_gp;               // emif_hps:emif_to_hps_gp -> agilex_hps:hps_emif_emif_to_gp
	wire  [4095:0] agilex_hps_hps_emif_hps_to_emif;            // agilex_hps:hps_emif_hps_to_emif -> emif_hps:hps_to_emif

	hps_sub_sys_agilex_axi_bridge_for_acp_0 agilex_axi_bridge_for_acp_0 (
		.clk             (acp_0_clock_clk),                         //   input,    width = 1,     clock.clk
		.reset           (acp_0_reset_reset),                       //   input,    width = 1,     reset.reset
		.csr_clk         (acp_0_csr_clock_clk),                     //   input,    width = 1, csr_clock.clk
		.csr_reset       (acp_0_csr_reset_reset),                   //   input,    width = 1, csr_reset.reset
		.addr            (acp_0_csr_address),                       //   input,    width = 1,       csr.address
		.read            (acp_0_csr_read),                          //   input,    width = 1,          .read
		.write           (acp_0_csr_write),                         //   input,    width = 1,          .write
		.writedata       (acp_0_csr_writedata),                     //   input,   width = 32,          .writedata
		.readdata        (acp_0_csr_readdata),                      //  output,   width = 32,          .readdata
		.axm_m0_araddr   (agilex_axi_bridge_for_acp_0_m0_araddr),   //  output,   width = 37,        m0.araddr
		.axm_m0_arburst  (agilex_axi_bridge_for_acp_0_m0_arburst),  //  output,    width = 2,          .arburst
		.axm_m0_arcache  (agilex_axi_bridge_for_acp_0_m0_arcache),  //  output,    width = 4,          .arcache
		.axm_m0_arid     (agilex_axi_bridge_for_acp_0_m0_arid),     //  output,    width = 5,          .arid
		.axm_m0_arlen    (agilex_axi_bridge_for_acp_0_m0_arlen),    //  output,    width = 8,          .arlen
		.axm_m0_arlock   (agilex_axi_bridge_for_acp_0_m0_arlock),   //  output,    width = 1,          .arlock
		.axm_m0_arprot   (agilex_axi_bridge_for_acp_0_m0_arprot),   //  output,    width = 3,          .arprot
		.axm_m0_arqos    (agilex_axi_bridge_for_acp_0_m0_arqos),    //  output,    width = 4,          .arqos
		.axm_m0_arready  (agilex_axi_bridge_for_acp_0_m0_arready),  //   input,    width = 1,          .arready
		.axm_m0_arsize   (agilex_axi_bridge_for_acp_0_m0_arsize),   //  output,    width = 3,          .arsize
		.axm_m0_arvalid  (agilex_axi_bridge_for_acp_0_m0_arvalid),  //  output,    width = 1,          .arvalid
		.axm_m0_arsnoop  (agilex_axi_bridge_for_acp_0_m0_arsnoop),  //  output,    width = 4,          .arsnoop
		.axm_m0_ardomain (agilex_axi_bridge_for_acp_0_m0_ardomain), //  output,    width = 2,          .ardomain
		.axm_m0_arbar    (agilex_axi_bridge_for_acp_0_m0_arbar),    //  output,    width = 2,          .arbar
		.axm_m0_aruser   (agilex_axi_bridge_for_acp_0_m0_aruser),   //  output,   width = 23,          .aruser
		.axm_m0_awaddr   (agilex_axi_bridge_for_acp_0_m0_awaddr),   //  output,   width = 37,          .awaddr
		.axm_m0_awburst  (agilex_axi_bridge_for_acp_0_m0_awburst),  //  output,    width = 2,          .awburst
		.axm_m0_awcache  (agilex_axi_bridge_for_acp_0_m0_awcache),  //  output,    width = 4,          .awcache
		.axm_m0_awid     (agilex_axi_bridge_for_acp_0_m0_awid),     //  output,    width = 5,          .awid
		.axm_m0_awlen    (agilex_axi_bridge_for_acp_0_m0_awlen),    //  output,    width = 8,          .awlen
		.axm_m0_awlock   (agilex_axi_bridge_for_acp_0_m0_awlock),   //  output,    width = 1,          .awlock
		.axm_m0_awprot   (agilex_axi_bridge_for_acp_0_m0_awprot),   //  output,    width = 3,          .awprot
		.axm_m0_awready  (agilex_axi_bridge_for_acp_0_m0_awready),  //   input,    width = 1,          .awready
		.axm_m0_awsize   (agilex_axi_bridge_for_acp_0_m0_awsize),   //  output,    width = 3,          .awsize
		.axm_m0_awvalid  (agilex_axi_bridge_for_acp_0_m0_awvalid),  //  output,    width = 1,          .awvalid
		.axm_m0_awqos    (agilex_axi_bridge_for_acp_0_m0_awqos),    //  output,    width = 4,          .awqos
		.axm_m0_bid      (agilex_axi_bridge_for_acp_0_m0_bid),      //   input,    width = 5,          .bid
		.axm_m0_bready   (agilex_axi_bridge_for_acp_0_m0_bready),   //  output,    width = 1,          .bready
		.axm_m0_bresp    (agilex_axi_bridge_for_acp_0_m0_bresp),    //   input,    width = 2,          .bresp
		.axm_m0_bvalid   (agilex_axi_bridge_for_acp_0_m0_bvalid),   //   input,    width = 1,          .bvalid
		.axm_m0_rdata    (agilex_axi_bridge_for_acp_0_m0_rdata),    //   input,  width = 512,          .rdata
		.axm_m0_rid      (agilex_axi_bridge_for_acp_0_m0_rid),      //   input,    width = 5,          .rid
		.axm_m0_rlast    (agilex_axi_bridge_for_acp_0_m0_rlast),    //   input,    width = 1,          .rlast
		.axm_m0_rready   (agilex_axi_bridge_for_acp_0_m0_rready),   //  output,    width = 1,          .rready
		.axm_m0_rresp    (agilex_axi_bridge_for_acp_0_m0_rresp),    //   input,    width = 2,          .rresp
		.axm_m0_rvalid   (agilex_axi_bridge_for_acp_0_m0_rvalid),   //   input,    width = 1,          .rvalid
		.axm_m0_wdata    (agilex_axi_bridge_for_acp_0_m0_wdata),    //  output,  width = 512,          .wdata
		.axm_m0_wlast    (agilex_axi_bridge_for_acp_0_m0_wlast),    //  output,    width = 1,          .wlast
		.axm_m0_wready   (agilex_axi_bridge_for_acp_0_m0_wready),   //   input,    width = 1,          .wready
		.axm_m0_wstrb    (agilex_axi_bridge_for_acp_0_m0_wstrb),    //  output,   width = 64,          .wstrb
		.axm_m0_wvalid   (agilex_axi_bridge_for_acp_0_m0_wvalid),   //  output,    width = 1,          .wvalid
		.axm_m0_awsnoop  (agilex_axi_bridge_for_acp_0_m0_awsnoop),  //  output,    width = 3,          .awsnoop
		.axm_m0_awdomain (agilex_axi_bridge_for_acp_0_m0_awdomain), //  output,    width = 2,          .awdomain
		.axm_m0_awbar    (agilex_axi_bridge_for_acp_0_m0_awbar),    //  output,    width = 2,          .awbar
		.axm_m0_awuser   (agilex_axi_bridge_for_acp_0_m0_awuser),   //  output,   width = 23,          .awuser
		.axs_s0_araddr   (acp_0_s0_araddr),                         //   input,   width = 37,        s0.araddr
		.axs_s0_arburst  (acp_0_s0_arburst),                        //   input,    width = 2,          .arburst
		.axs_s0_arcache  (acp_0_s0_arcache),                        //   input,    width = 4,          .arcache
		.axs_s0_arid     (acp_0_s0_arid),                           //   input,    width = 4,          .arid
		.axs_s0_arlen    (acp_0_s0_arlen),                          //   input,    width = 8,          .arlen
		.axs_s0_arlock   (acp_0_s0_arlock),                         //   input,    width = 1,          .arlock
		.axs_s0_arprot   (acp_0_s0_arprot),                         //   input,    width = 3,          .arprot
		.axs_s0_arready  (acp_0_s0_arready),                        //  output,    width = 1,          .arready
		.axs_s0_arsize   (acp_0_s0_arsize),                         //   input,    width = 3,          .arsize
		.axs_s0_arvalid  (acp_0_s0_arvalid),                        //   input,    width = 1,          .arvalid
		.axs_s0_awaddr   (acp_0_s0_awaddr),                         //   input,   width = 37,          .awaddr
		.axs_s0_awburst  (acp_0_s0_awburst),                        //   input,    width = 2,          .awburst
		.axs_s0_awcache  (acp_0_s0_awcache),                        //   input,    width = 4,          .awcache
		.axs_s0_awid     (acp_0_s0_awid),                           //   input,    width = 4,          .awid
		.axs_s0_awlen    (acp_0_s0_awlen),                          //   input,    width = 8,          .awlen
		.axs_s0_awlock   (acp_0_s0_awlock),                         //   input,    width = 1,          .awlock
		.axs_s0_awprot   (acp_0_s0_awprot),                         //   input,    width = 3,          .awprot
		.axs_s0_awready  (acp_0_s0_awready),                        //  output,    width = 1,          .awready
		.axs_s0_awsize   (acp_0_s0_awsize),                         //   input,    width = 3,          .awsize
		.axs_s0_awvalid  (acp_0_s0_awvalid),                        //   input,    width = 1,          .awvalid
		.axs_s0_bid      (acp_0_s0_bid),                            //  output,    width = 4,          .bid
		.axs_s0_bready   (acp_0_s0_bready),                         //   input,    width = 1,          .bready
		.axs_s0_bresp    (acp_0_s0_bresp),                          //  output,    width = 2,          .bresp
		.axs_s0_bvalid   (acp_0_s0_bvalid),                         //  output,    width = 1,          .bvalid
		.axs_s0_rdata    (acp_0_s0_rdata),                          //  output,  width = 512,          .rdata
		.axs_s0_rid      (acp_0_s0_rid),                            //  output,    width = 4,          .rid
		.axs_s0_rlast    (acp_0_s0_rlast),                          //  output,    width = 1,          .rlast
		.axs_s0_rready   (acp_0_s0_rready),                         //   input,    width = 1,          .rready
		.axs_s0_rresp    (acp_0_s0_rresp),                          //  output,    width = 2,          .rresp
		.axs_s0_rvalid   (acp_0_s0_rvalid),                         //  output,    width = 1,          .rvalid
		.axs_s0_wdata    (acp_0_s0_wdata),                          //   input,  width = 512,          .wdata
		.axs_s0_wlast    (acp_0_s0_wlast),                          //   input,    width = 1,          .wlast
		.axs_s0_wready   (acp_0_s0_wready),                         //  output,    width = 1,          .wready
		.axs_s0_wstrb    (acp_0_s0_wstrb),                          //   input,   width = 64,          .wstrb
		.axs_s0_wvalid   (acp_0_s0_wvalid)                          //   input,    width = 1,          .wvalid
	);

	agilex_hps agilex_hps (
		.s2f_user_clk0_hio       (),                                          //  output,     width = 1,   h2f_user0_clock.clk
		.s2f_user_clk1_hio       (),                                          //  output,     width = 1,   h2f_user1_clock.clk
		.h2f_mpu_fpga_eventi     (),                                          //   input,     width = 1,    h2f_mpu_events.fpga_eventi
		.h2f_mpu_fpga_evento     (),                                          //  output,     width = 1,                  .fpga_evento
		.h2f_mpu_fpga_standbywfe (),                                          //  output,     width = 4,                  .fpga_standbywfe
		.h2f_mpu_fpga_standbywfi (),                                          //  output,     width = 4,                  .fpga_standbywfi
		.f2h_stm_hwevents        (agilex_hps_f2h_stm_hw_events_stm_hwevents), //   input,    width = 44, f2h_stm_hw_events.stm_hwevents
		.h2f_cs_ntrst            (agilex_hps_h2f_cs_ntrst),                   //   input,     width = 1,            h2f_cs.ntrst
		.h2f_cs_tck              (agilex_hps_h2f_cs_tck),                     //   input,     width = 1,                  .tck
		.h2f_cs_tdi              (agilex_hps_h2f_cs_tdi),                     //   input,     width = 1,                  .tdi
		.h2f_cs_tdo              (agilex_hps_h2f_cs_tdo),                     //  output,     width = 1,                  .tdo
		.h2f_cs_tdoen            (agilex_hps_h2f_cs_tdoen),                   //  output,     width = 1,                  .tdoen
		.h2f_cs_tms              (agilex_hps_h2f_cs_tms),                     //   input,     width = 1,                  .tms
		.hps_emif_emif_to_hps    (emif_hps_hps_emif_emif_to_hps),             //   input,  width = 4096,          hps_emif.emif_to_hps
		.hps_emif_hps_to_emif    (agilex_hps_hps_emif_hps_to_emif),           //  output,  width = 4096,                  .hps_to_emif
		.hps_emif_emif_to_gp     (emif_hps_hps_emif_emif_to_gp),              //   input,     width = 1,                  .emif_to_gp
		.hps_emif_gp_to_emif     (agilex_hps_hps_emif_gp_to_emif),            //  output,     width = 2,                  .gp_to_emif
		.EMAC1_TX_CLK            (agilex_hps_hps_io_EMAC1_TX_CLK),            //  output,     width = 1,            hps_io.EMAC1_TX_CLK
		.EMAC1_TXD0              (agilex_hps_hps_io_EMAC1_TXD0),              //  output,     width = 1,                  .EMAC1_TXD0
		.EMAC1_TXD1              (agilex_hps_hps_io_EMAC1_TXD1),              //  output,     width = 1,                  .EMAC1_TXD1
		.EMAC1_TXD2              (agilex_hps_hps_io_EMAC1_TXD2),              //  output,     width = 1,                  .EMAC1_TXD2
		.EMAC1_TXD3              (agilex_hps_hps_io_EMAC1_TXD3),              //  output,     width = 1,                  .EMAC1_TXD3
		.EMAC1_RX_CTL            (agilex_hps_hps_io_EMAC1_RX_CTL),            //   input,     width = 1,                  .EMAC1_RX_CTL
		.EMAC1_TX_CTL            (agilex_hps_hps_io_EMAC1_TX_CTL),            //  output,     width = 1,                  .EMAC1_TX_CTL
		.EMAC1_RX_CLK            (agilex_hps_hps_io_EMAC1_RX_CLK),            //   input,     width = 1,                  .EMAC1_RX_CLK
		.EMAC1_RXD0              (agilex_hps_hps_io_EMAC1_RXD0),              //   input,     width = 1,                  .EMAC1_RXD0
		.EMAC1_RXD1              (agilex_hps_hps_io_EMAC1_RXD1),              //   input,     width = 1,                  .EMAC1_RXD1
		.EMAC1_RXD2              (agilex_hps_hps_io_EMAC1_RXD2),              //   input,     width = 1,                  .EMAC1_RXD2
		.EMAC1_RXD3              (agilex_hps_hps_io_EMAC1_RXD3),              //   input,     width = 1,                  .EMAC1_RXD3
		.EMAC1_MDIO              (agilex_hps_hps_io_EMAC1_MDIO),              //   inout,     width = 1,                  .EMAC1_MDIO
		.EMAC1_MDC               (agilex_hps_hps_io_EMAC1_MDC),               //  output,     width = 1,                  .EMAC1_MDC
		.SDMMC_CMD               (agilex_hps_hps_io_SDMMC_CMD),               //   inout,     width = 1,                  .SDMMC_CMD
		.SDMMC_D0                (agilex_hps_hps_io_SDMMC_D0),                //   inout,     width = 1,                  .SDMMC_D0
		.SDMMC_D1                (agilex_hps_hps_io_SDMMC_D1),                //   inout,     width = 1,                  .SDMMC_D1
		.SDMMC_D2                (agilex_hps_hps_io_SDMMC_D2),                //   inout,     width = 1,                  .SDMMC_D2
		.SDMMC_D3                (agilex_hps_hps_io_SDMMC_D3),                //   inout,     width = 1,                  .SDMMC_D3
		.SDMMC_D4                (agilex_hps_hps_io_SDMMC_D4),                //   inout,     width = 1,                  .SDMMC_D4
		.SDMMC_D5                (agilex_hps_hps_io_SDMMC_D5),                //   inout,     width = 1,                  .SDMMC_D5
		.SDMMC_D6                (agilex_hps_hps_io_SDMMC_D6),                //   inout,     width = 1,                  .SDMMC_D6
		.SDMMC_D7                (agilex_hps_hps_io_SDMMC_D7),                //   inout,     width = 1,                  .SDMMC_D7
		.SDMMC_CCLK              (agilex_hps_hps_io_SDMMC_CCLK),              //  output,     width = 1,                  .SDMMC_CCLK
		.SPIM0_CLK               (agilex_hps_hps_io_SPIM0_CLK),               //  output,     width = 1,                  .SPIM0_CLK
		.SPIM0_MOSI              (agilex_hps_hps_io_SPIM0_MOSI),              //  output,     width = 1,                  .SPIM0_MOSI
		.SPIM0_MISO              (agilex_hps_hps_io_SPIM0_MISO),              //   input,     width = 1,                  .SPIM0_MISO
		.SPIM0_SS0_N             (agilex_hps_hps_io_SPIM0_SS0_N),             //  output,     width = 1,                  .SPIM0_SS0_N
		.SPIM1_CLK               (agilex_hps_hps_io_SPIM1_CLK),               //  output,     width = 1,                  .SPIM1_CLK
		.SPIM1_MOSI              (agilex_hps_hps_io_SPIM1_MOSI),              //  output,     width = 1,                  .SPIM1_MOSI
		.SPIM1_MISO              (agilex_hps_hps_io_SPIM1_MISO),              //   input,     width = 1,                  .SPIM1_MISO
		.SPIM1_SS0_N             (agilex_hps_hps_io_SPIM1_SS0_N),             //  output,     width = 1,                  .SPIM1_SS0_N
		.SPIM1_SS1_N             (agilex_hps_hps_io_SPIM1_SS1_N),             //  output,     width = 1,                  .SPIM1_SS1_N
		.UART1_RX                (agilex_hps_hps_io_UART1_RX),                //   input,     width = 1,                  .UART1_RX
		.UART1_TX                (agilex_hps_hps_io_UART1_TX),                //  output,     width = 1,                  .UART1_TX
		.I2C1_SDA                (agilex_hps_hps_io_I2C1_SDA),                //   inout,     width = 1,                  .I2C1_SDA
		.I2C1_SCL                (agilex_hps_hps_io_I2C1_SCL),                //   inout,     width = 1,                  .I2C1_SCL
		.hps_osc_clk             (agilex_hps_hps_io_hps_osc_clk),             //   input,     width = 1,                  .hps_osc_clk
		.gpio0_io11              (agilex_hps_hps_io_gpio0_io11),              //   inout,     width = 1,                  .gpio0_io11
		.gpio0_io12              (agilex_hps_hps_io_gpio0_io12),              //   inout,     width = 1,                  .gpio0_io12
		.gpio0_io13              (agilex_hps_hps_io_gpio0_io13),              //   inout,     width = 1,                  .gpio0_io13
		.gpio0_io14              (agilex_hps_hps_io_gpio0_io14),              //   inout,     width = 1,                  .gpio0_io14
		.gpio0_io15              (agilex_hps_hps_io_gpio0_io15),              //   inout,     width = 1,                  .gpio0_io15
		.gpio0_io16              (agilex_hps_hps_io_gpio0_io16),              //   inout,     width = 1,                  .gpio0_io16
		.gpio0_io17              (agilex_hps_hps_io_gpio0_io17),              //   inout,     width = 1,                  .gpio0_io17
		.gpio0_io18              (agilex_hps_hps_io_gpio0_io18),              //   inout,     width = 1,                  .gpio0_io18
		.gpio1_io16              (agilex_hps_hps_io_gpio1_io16),              //   inout,     width = 1,                  .gpio1_io16
		.gpio1_io17              (agilex_hps_hps_io_gpio1_io17),              //   inout,     width = 1,                  .gpio1_io17
		.h2f_rst                 (agilex_hps_h2f_reset_reset),                //  output,     width = 1,         h2f_reset.reset
		.h2f_axi_clk             (agilex_hps_h2f_axi_clock_clk),              //   input,     width = 1,     h2f_axi_clock.clk
		.h2f_axi_rst_n           (agilex_hps_h2f_axi_reset_reset_n),          //   input,     width = 1,     h2f_axi_reset.reset_n
		.h2f_AWID                (agilex_hps_h2f_axi_master_awid),            //  output,     width = 4,    h2f_axi_master.awid
		.h2f_AWADDR              (agilex_hps_h2f_axi_master_awaddr),          //  output,    width = 32,                  .awaddr
		.h2f_AWLEN               (agilex_hps_h2f_axi_master_awlen),           //  output,     width = 8,                  .awlen
		.h2f_AWSIZE              (agilex_hps_h2f_axi_master_awsize),          //  output,     width = 3,                  .awsize
		.h2f_AWBURST             (agilex_hps_h2f_axi_master_awburst),         //  output,     width = 2,                  .awburst
		.h2f_AWLOCK              (agilex_hps_h2f_axi_master_awlock),          //  output,     width = 1,                  .awlock
		.h2f_AWCACHE             (agilex_hps_h2f_axi_master_awcache),         //  output,     width = 4,                  .awcache
		.h2f_AWPROT              (agilex_hps_h2f_axi_master_awprot),          //  output,     width = 3,                  .awprot
		.h2f_AWVALID             (agilex_hps_h2f_axi_master_awvalid),         //  output,     width = 1,                  .awvalid
		.h2f_AWREADY             (agilex_hps_h2f_axi_master_awready),         //   input,     width = 1,                  .awready
		.h2f_WDATA               (agilex_hps_h2f_axi_master_wdata),           //  output,   width = 128,                  .wdata
		.h2f_WSTRB               (agilex_hps_h2f_axi_master_wstrb),           //  output,    width = 16,                  .wstrb
		.h2f_WLAST               (agilex_hps_h2f_axi_master_wlast),           //  output,     width = 1,                  .wlast
		.h2f_WVALID              (agilex_hps_h2f_axi_master_wvalid),          //  output,     width = 1,                  .wvalid
		.h2f_WREADY              (agilex_hps_h2f_axi_master_wready),          //   input,     width = 1,                  .wready
		.h2f_BID                 (agilex_hps_h2f_axi_master_bid),             //   input,     width = 4,                  .bid
		.h2f_BRESP               (agilex_hps_h2f_axi_master_bresp),           //   input,     width = 2,                  .bresp
		.h2f_BVALID              (agilex_hps_h2f_axi_master_bvalid),          //   input,     width = 1,                  .bvalid
		.h2f_BREADY              (agilex_hps_h2f_axi_master_bready),          //  output,     width = 1,                  .bready
		.h2f_ARID                (agilex_hps_h2f_axi_master_arid),            //  output,     width = 4,                  .arid
		.h2f_ARADDR              (agilex_hps_h2f_axi_master_araddr),          //  output,    width = 32,                  .araddr
		.h2f_ARLEN               (agilex_hps_h2f_axi_master_arlen),           //  output,     width = 8,                  .arlen
		.h2f_ARSIZE              (agilex_hps_h2f_axi_master_arsize),          //  output,     width = 3,                  .arsize
		.h2f_ARBURST             (agilex_hps_h2f_axi_master_arburst),         //  output,     width = 2,                  .arburst
		.h2f_ARLOCK              (agilex_hps_h2f_axi_master_arlock),          //  output,     width = 1,                  .arlock
		.h2f_ARCACHE             (agilex_hps_h2f_axi_master_arcache),         //  output,     width = 4,                  .arcache
		.h2f_ARPROT              (agilex_hps_h2f_axi_master_arprot),          //  output,     width = 3,                  .arprot
		.h2f_ARVALID             (agilex_hps_h2f_axi_master_arvalid),         //  output,     width = 1,                  .arvalid
		.h2f_ARREADY             (agilex_hps_h2f_axi_master_arready),         //   input,     width = 1,                  .arready
		.h2f_RID                 (agilex_hps_h2f_axi_master_rid),             //   input,     width = 4,                  .rid
		.h2f_RDATA               (agilex_hps_h2f_axi_master_rdata),           //   input,   width = 128,                  .rdata
		.h2f_RRESP               (agilex_hps_h2f_axi_master_rresp),           //   input,     width = 2,                  .rresp
		.h2f_RLAST               (agilex_hps_h2f_axi_master_rlast),           //   input,     width = 1,                  .rlast
		.h2f_RVALID              (agilex_hps_h2f_axi_master_rvalid),          //   input,     width = 1,                  .rvalid
		.h2f_RREADY              (agilex_hps_h2f_axi_master_rready),          //  output,     width = 1,                  .rready
		.h2f_lw_axi_clk          (agilex_hps_h2f_lw_axi_clock_clk),           //   input,     width = 1,  h2f_lw_axi_clock.clk
		.h2f_lw_axi_rst_n        (agilex_hps_h2f_lw_axi_reset_reset_n),       //   input,     width = 1,  h2f_lw_axi_reset.reset_n
		.h2f_lw_AWID             (agilex_hps_h2f_lw_axi_master_awid),         //  output,     width = 4, h2f_lw_axi_master.awid
		.h2f_lw_AWADDR           (agilex_hps_h2f_lw_axi_master_awaddr),       //  output,    width = 21,                  .awaddr
		.h2f_lw_AWLEN            (agilex_hps_h2f_lw_axi_master_awlen),        //  output,     width = 8,                  .awlen
		.h2f_lw_AWSIZE           (agilex_hps_h2f_lw_axi_master_awsize),       //  output,     width = 3,                  .awsize
		.h2f_lw_AWBURST          (agilex_hps_h2f_lw_axi_master_awburst),      //  output,     width = 2,                  .awburst
		.h2f_lw_AWLOCK           (agilex_hps_h2f_lw_axi_master_awlock),       //  output,     width = 1,                  .awlock
		.h2f_lw_AWCACHE          (agilex_hps_h2f_lw_axi_master_awcache),      //  output,     width = 4,                  .awcache
		.h2f_lw_AWPROT           (agilex_hps_h2f_lw_axi_master_awprot),       //  output,     width = 3,                  .awprot
		.h2f_lw_AWVALID          (agilex_hps_h2f_lw_axi_master_awvalid),      //  output,     width = 1,                  .awvalid
		.h2f_lw_AWREADY          (agilex_hps_h2f_lw_axi_master_awready),      //   input,     width = 1,                  .awready
		.h2f_lw_WDATA            (agilex_hps_h2f_lw_axi_master_wdata),        //  output,    width = 32,                  .wdata
		.h2f_lw_WSTRB            (agilex_hps_h2f_lw_axi_master_wstrb),        //  output,     width = 4,                  .wstrb
		.h2f_lw_WLAST            (agilex_hps_h2f_lw_axi_master_wlast),        //  output,     width = 1,                  .wlast
		.h2f_lw_WVALID           (agilex_hps_h2f_lw_axi_master_wvalid),       //  output,     width = 1,                  .wvalid
		.h2f_lw_WREADY           (agilex_hps_h2f_lw_axi_master_wready),       //   input,     width = 1,                  .wready
		.h2f_lw_BID              (agilex_hps_h2f_lw_axi_master_bid),          //   input,     width = 4,                  .bid
		.h2f_lw_BRESP            (agilex_hps_h2f_lw_axi_master_bresp),        //   input,     width = 2,                  .bresp
		.h2f_lw_BVALID           (agilex_hps_h2f_lw_axi_master_bvalid),       //   input,     width = 1,                  .bvalid
		.h2f_lw_BREADY           (agilex_hps_h2f_lw_axi_master_bready),       //  output,     width = 1,                  .bready
		.h2f_lw_ARID             (agilex_hps_h2f_lw_axi_master_arid),         //  output,     width = 4,                  .arid
		.h2f_lw_ARADDR           (agilex_hps_h2f_lw_axi_master_araddr),       //  output,    width = 21,                  .araddr
		.h2f_lw_ARLEN            (agilex_hps_h2f_lw_axi_master_arlen),        //  output,     width = 8,                  .arlen
		.h2f_lw_ARSIZE           (agilex_hps_h2f_lw_axi_master_arsize),       //  output,     width = 3,                  .arsize
		.h2f_lw_ARBURST          (agilex_hps_h2f_lw_axi_master_arburst),      //  output,     width = 2,                  .arburst
		.h2f_lw_ARLOCK           (agilex_hps_h2f_lw_axi_master_arlock),       //  output,     width = 1,                  .arlock
		.h2f_lw_ARCACHE          (agilex_hps_h2f_lw_axi_master_arcache),      //  output,     width = 4,                  .arcache
		.h2f_lw_ARPROT           (agilex_hps_h2f_lw_axi_master_arprot),       //  output,     width = 3,                  .arprot
		.h2f_lw_ARVALID          (agilex_hps_h2f_lw_axi_master_arvalid),      //  output,     width = 1,                  .arvalid
		.h2f_lw_ARREADY          (agilex_hps_h2f_lw_axi_master_arready),      //   input,     width = 1,                  .arready
		.h2f_lw_RID              (agilex_hps_h2f_lw_axi_master_rid),          //   input,     width = 4,                  .rid
		.h2f_lw_RDATA            (agilex_hps_h2f_lw_axi_master_rdata),        //   input,    width = 32,                  .rdata
		.h2f_lw_RRESP            (agilex_hps_h2f_lw_axi_master_rresp),        //   input,     width = 2,                  .rresp
		.h2f_lw_RLAST            (agilex_hps_h2f_lw_axi_master_rlast),        //   input,     width = 1,                  .rlast
		.h2f_lw_RVALID           (agilex_hps_h2f_lw_axi_master_rvalid),       //   input,     width = 1,                  .rvalid
		.h2f_lw_RREADY           (agilex_hps_h2f_lw_axi_master_rready),       //  output,     width = 1,                  .rready
		.f2h_axi_clk             (agilex_hps_f2h_axi_clock_clk),              //   input,     width = 1,     f2h_axi_clock.clk
		.f2h_axi_rst_n           (agilex_hps_f2h_axi_reset_reset_n),          //   input,     width = 1,     f2h_axi_reset.reset_n
		.f2h_AWID                (agilex_axi_bridge_for_acp_0_m0_awid),       //   input,     width = 5,     f2h_axi_slave.awid
		.f2h_AWADDR              (agilex_axi_bridge_for_acp_0_m0_awaddr),     //   input,    width = 37,                  .awaddr
		.f2h_AWLEN               (agilex_axi_bridge_for_acp_0_m0_awlen),      //   input,     width = 8,                  .awlen
		.f2h_AWSIZE              (agilex_axi_bridge_for_acp_0_m0_awsize),     //   input,     width = 3,                  .awsize
		.f2h_AWBURST             (agilex_axi_bridge_for_acp_0_m0_awburst),    //   input,     width = 2,                  .awburst
		.f2h_AWLOCK              (agilex_axi_bridge_for_acp_0_m0_awlock),     //   input,     width = 1,                  .awlock
		.f2h_AWCACHE             (agilex_axi_bridge_for_acp_0_m0_awcache),    //   input,     width = 4,                  .awcache
		.f2h_AWPROT              (agilex_axi_bridge_for_acp_0_m0_awprot),     //   input,     width = 3,                  .awprot
		.f2h_AWVALID             (agilex_axi_bridge_for_acp_0_m0_awvalid),    //   input,     width = 1,                  .awvalid
		.f2h_AWREADY             (agilex_axi_bridge_for_acp_0_m0_awready),    //  output,     width = 1,                  .awready
		.f2h_AWQOS               (agilex_axi_bridge_for_acp_0_m0_awqos),      //   input,     width = 4,                  .awqos
		.f2h_WDATA               (agilex_axi_bridge_for_acp_0_m0_wdata),      //   input,   width = 512,                  .wdata
		.f2h_WSTRB               (agilex_axi_bridge_for_acp_0_m0_wstrb),      //   input,    width = 64,                  .wstrb
		.f2h_WLAST               (agilex_axi_bridge_for_acp_0_m0_wlast),      //   input,     width = 1,                  .wlast
		.f2h_WVALID              (agilex_axi_bridge_for_acp_0_m0_wvalid),     //   input,     width = 1,                  .wvalid
		.f2h_WREADY              (agilex_axi_bridge_for_acp_0_m0_wready),     //  output,     width = 1,                  .wready
		.f2h_BID                 (agilex_axi_bridge_for_acp_0_m0_bid),        //  output,     width = 5,                  .bid
		.f2h_BRESP               (agilex_axi_bridge_for_acp_0_m0_bresp),      //  output,     width = 2,                  .bresp
		.f2h_BVALID              (agilex_axi_bridge_for_acp_0_m0_bvalid),     //  output,     width = 1,                  .bvalid
		.f2h_BREADY              (agilex_axi_bridge_for_acp_0_m0_bready),     //   input,     width = 1,                  .bready
		.f2h_ARID                (agilex_axi_bridge_for_acp_0_m0_arid),       //   input,     width = 5,                  .arid
		.f2h_ARADDR              (agilex_axi_bridge_for_acp_0_m0_araddr),     //   input,    width = 37,                  .araddr
		.f2h_ARLEN               (agilex_axi_bridge_for_acp_0_m0_arlen),      //   input,     width = 8,                  .arlen
		.f2h_ARSIZE              (agilex_axi_bridge_for_acp_0_m0_arsize),     //   input,     width = 3,                  .arsize
		.f2h_ARBURST             (agilex_axi_bridge_for_acp_0_m0_arburst),    //   input,     width = 2,                  .arburst
		.f2h_ARLOCK              (agilex_axi_bridge_for_acp_0_m0_arlock),     //   input,     width = 1,                  .arlock
		.f2h_ARCACHE             (agilex_axi_bridge_for_acp_0_m0_arcache),    //   input,     width = 4,                  .arcache
		.f2h_ARPROT              (agilex_axi_bridge_for_acp_0_m0_arprot),     //   input,     width = 3,                  .arprot
		.f2h_ARVALID             (agilex_axi_bridge_for_acp_0_m0_arvalid),    //   input,     width = 1,                  .arvalid
		.f2h_ARREADY             (agilex_axi_bridge_for_acp_0_m0_arready),    //  output,     width = 1,                  .arready
		.f2h_ARQOS               (agilex_axi_bridge_for_acp_0_m0_arqos),      //   input,     width = 4,                  .arqos
		.f2h_RID                 (agilex_axi_bridge_for_acp_0_m0_rid),        //  output,     width = 5,                  .rid
		.f2h_RDATA               (agilex_axi_bridge_for_acp_0_m0_rdata),      //  output,   width = 512,                  .rdata
		.f2h_RRESP               (agilex_axi_bridge_for_acp_0_m0_rresp),      //  output,     width = 2,                  .rresp
		.f2h_RLAST               (agilex_axi_bridge_for_acp_0_m0_rlast),      //  output,     width = 1,                  .rlast
		.f2h_RVALID              (agilex_axi_bridge_for_acp_0_m0_rvalid),     //  output,     width = 1,                  .rvalid
		.f2h_RREADY              (agilex_axi_bridge_for_acp_0_m0_rready),     //   input,     width = 1,                  .rready
		.f2h_AWDOMAIN            (agilex_axi_bridge_for_acp_0_m0_awdomain),   //   input,     width = 2,                  .awdomain
		.f2h_AWBAR               (agilex_axi_bridge_for_acp_0_m0_awbar),      //   input,     width = 2,                  .awbar
		.f2h_ARDOMAIN            (agilex_axi_bridge_for_acp_0_m0_ardomain),   //   input,     width = 2,                  .ardomain
		.f2h_ARBAR               (agilex_axi_bridge_for_acp_0_m0_arbar),      //   input,     width = 2,                  .arbar
		.f2h_ARSNOOP             (agilex_axi_bridge_for_acp_0_m0_arsnoop),    //   input,     width = 4,                  .arsnoop
		.f2h_AWSNOOP             (agilex_axi_bridge_for_acp_0_m0_awsnoop),    //   input,     width = 3,                  .awsnoop
		.f2h_ARUSER              (agilex_axi_bridge_for_acp_0_m0_aruser),     //   input,    width = 23,                  .aruser
		.f2h_AWUSER              (agilex_axi_bridge_for_acp_0_m0_awuser),     //   input,    width = 23,                  .awuser
		.f2h_irq_p0              (agilex_hps_f2h_irq0_irq),                   //   input,    width = 32,          f2h_irq0.irq
		.f2h_irq_p1              (agilex_hps_f2h_irq1_irq)                    //   input,    width = 32,          f2h_irq1.irq
	);

	emif_calbus_0 emif_calbus_0 (
		.calbus_read_0          (emif_calbus_0_emif_calbus_0_calbus_read),    //  output,     width = 1,   emif_calbus_0.calbus_read
		.calbus_write_0         (emif_calbus_0_emif_calbus_0_calbus_write),   //  output,     width = 1,                .calbus_write
		.calbus_address_0       (emif_calbus_0_emif_calbus_0_calbus_address), //  output,    width = 20,                .calbus_address
		.calbus_wdata_0         (emif_calbus_0_emif_calbus_0_calbus_wdata),   //  output,    width = 32,                .calbus_wdata
		.calbus_rdata_0         (emif_hps_emif_calbus_calbus_rdata),          //   input,    width = 32,                .calbus_rdata
		.calbus_seq_param_tbl_0 (emif_hps_emif_calbus_calbus_seq_param_tbl),  //   input,  width = 4096,                .calbus_seq_param_tbl
		.calbus_clk             (emif_calbus_0_emif_calbus_clk_clk)           //  output,     width = 1, emif_calbus_clk.clk
	);

	emif_hps emif_hps (
		.pll_ref_clk          (emif_hps_pll_ref_clk_clk),                   //   input,     width = 1,     pll_ref_clk.clk
		.oct_rzqin            (emif_hps_oct_oct_rzqin),                     //   input,     width = 1,             oct.oct_rzqin
		.mem_ck               (emif_hps_mem_mem_ck),                        //  output,     width = 1,             mem.mem_ck
		.mem_ck_n             (emif_hps_mem_mem_ck_n),                      //  output,     width = 1,                .mem_ck_n
		.mem_a                (emif_hps_mem_mem_a),                         //  output,    width = 17,                .mem_a
		.mem_act_n            (emif_hps_mem_mem_act_n),                     //  output,     width = 1,                .mem_act_n
		.mem_ba               (emif_hps_mem_mem_ba),                        //  output,     width = 2,                .mem_ba
		.mem_bg               (emif_hps_mem_mem_bg),                        //  output,     width = 1,                .mem_bg
		.mem_cke              (emif_hps_mem_mem_cke),                       //  output,     width = 1,                .mem_cke
		.mem_cs_n             (emif_hps_mem_mem_cs_n),                      //  output,     width = 2,                .mem_cs_n
		.mem_odt              (emif_hps_mem_mem_odt),                       //  output,     width = 1,                .mem_odt
		.mem_reset_n          (emif_hps_mem_mem_reset_n),                   //  output,     width = 1,                .mem_reset_n
		.mem_par              (emif_hps_mem_mem_par),                       //  output,     width = 1,                .mem_par
		.mem_alert_n          (emif_hps_mem_mem_alert_n),                   //   input,     width = 1,                .mem_alert_n
		.mem_dqs              (emif_hps_mem_mem_dqs),                       //   inout,     width = 9,                .mem_dqs
		.mem_dqs_n            (emif_hps_mem_mem_dqs_n),                     //   inout,     width = 9,                .mem_dqs_n
		.mem_dq               (emif_hps_mem_mem_dq),                        //   inout,    width = 72,                .mem_dq
		.mem_dbi_n            (emif_hps_mem_mem_dbi_n),                     //   inout,     width = 9,                .mem_dbi_n
		.hps_to_emif          (agilex_hps_hps_emif_hps_to_emif),            //   input,  width = 4096,        hps_emif.hps_to_emif
		.emif_to_hps          (emif_hps_hps_emif_emif_to_hps),              //  output,  width = 4096,                .emif_to_hps
		.hps_to_emif_gp       (agilex_hps_hps_emif_gp_to_emif),             //   input,     width = 2,                .gp_to_emif
		.emif_to_hps_gp       (emif_hps_hps_emif_emif_to_gp),               //  output,     width = 1,                .emif_to_gp
		.calbus_read          (emif_calbus_0_emif_calbus_0_calbus_read),    //   input,     width = 1,     emif_calbus.calbus_read
		.calbus_write         (emif_calbus_0_emif_calbus_0_calbus_write),   //   input,     width = 1,                .calbus_write
		.calbus_address       (emif_calbus_0_emif_calbus_0_calbus_address), //   input,    width = 20,                .calbus_address
		.calbus_wdata         (emif_calbus_0_emif_calbus_0_calbus_wdata),   //   input,    width = 32,                .calbus_wdata
		.calbus_rdata         (emif_hps_emif_calbus_calbus_rdata),          //  output,    width = 32,                .calbus_rdata
		.calbus_seq_param_tbl (emif_hps_emif_calbus_calbus_seq_param_tbl),  //  output,  width = 4096,                .calbus_seq_param_tbl
		.calbus_clk           (emif_calbus_0_emif_calbus_clk_clk)           //   input,     width = 1, emif_calbus_clk.clk
	);

endmodule
