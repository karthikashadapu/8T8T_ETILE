// sys_manager.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module sys_manager (
		input  wire        clk_100_in_clk_clk,                               //                           clk_100_in_clk.clk
		output wire        clk_100_out_clk_clk,                              //                          clk_100_out_clk.clk
		input  wire        dma_subsys_port0_rx_dma_resetn_clk_clk,           //       dma_subsys_port0_rx_dma_resetn_clk.clk
		input  wire        dma_subsys_port0_rx_dma_resetn_in_reset_reset_n,  //  dma_subsys_port0_rx_dma_resetn_in_reset.reset_n
		output wire        dma_subsys_port0_rx_dma_resetn_out_reset_reset_n, // dma_subsys_port0_rx_dma_resetn_out_reset.reset_n
		input  wire        dma_subsys_port1_rx_dma_resetn_clk_clk,           //       dma_subsys_port1_rx_dma_resetn_clk.clk
		input  wire        dma_subsys_port1_rx_dma_resetn_in_reset_reset_n,  //  dma_subsys_port1_rx_dma_resetn_in_reset.reset_n
		output wire        dma_subsys_port1_rx_dma_resetn_out_reset_reset_n, // dma_subsys_port1_rx_dma_resetn_out_reset.reset_n
		input  wire        ftile_iopll_ptp_sampling_refclk_clk,              //          ftile_iopll_ptp_sampling_refclk.clk
		input  wire        ftile_iopll_ptp_sampling_reset_reset,             //           ftile_iopll_ptp_sampling_reset.reset
		output wire        ftile_iopll_ptp_sampling_outclk0_clk,             //         ftile_iopll_ptp_sampling_outclk0.clk
		input  wire        ftile_iopll_todsync_sampling_refclk_clk,          //      ftile_iopll_todsync_sampling_refclk.clk
		output wire        ftile_iopll_todsync_sampling_locked_lock,         //      ftile_iopll_todsync_sampling_locked.lock
		input  wire        ftile_iopll_todsync_sampling_reset_reset,         //       ftile_iopll_todsync_sampling_reset.reset
		output wire        ftile_iopll_todsync_sampling_outclk0_clk,         //     ftile_iopll_todsync_sampling_outclk0.clk
		input  wire        qsys_top_master_todclk_0_in_clk_clk,              //          qsys_top_master_todclk_0_in_clk.clk
		output wire        qsys_top_master_todclk_0_out_clk_clk,             //         qsys_top_master_todclk_0_out_clk.clk
		input  wire        rst_in_clk_clk,                                   //                               rst_in_clk.clk
		input  wire        rst_in_in_reset_reset_n,                          //                          rst_in_in_reset.reset_n
		output wire        rst_in_out_reset_reset_n,                         //                         rst_in_out_reset.reset_n
		input  wire        sysid_clk_clk,                                    //                                sysid_clk.clk
		input  wire        sysid_reset_reset_n,                              //                              sysid_reset.reset_n
		output wire [31:0] sysid_control_slave_readdata,                     //                      sysid_control_slave.readdata
		input  wire        sysid_control_slave_address,                      //                                         .address
		output wire        user_rst_clkgate_0_ninit_done_ninit_done          //            user_rst_clkgate_0_ninit_done.ninit_done
	);

	clk_100 clk_100 (
		.in_clk  (clk_100_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (clk_100_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	dma_subsys_port0_rx_dma_resetn dma_subsys_port0_rx_dma_resetn (
		.clk         (dma_subsys_port0_rx_dma_resetn_clk_clk),           //   input,  width = 1,       clk.clk
		.in_reset_n  (dma_subsys_port0_rx_dma_resetn_in_reset_reset_n),  //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (dma_subsys_port0_rx_dma_resetn_out_reset_reset_n)  //  output,  width = 1, out_reset.reset_n
	);

	dma_subsys_port1_rx_dma_resetn dma_subsys_port1_rx_dma_resetn (
		.clk         (dma_subsys_port1_rx_dma_resetn_clk_clk),           //   input,  width = 1,       clk.clk
		.in_reset_n  (dma_subsys_port1_rx_dma_resetn_in_reset_reset_n),  //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (dma_subsys_port1_rx_dma_resetn_out_reset_reset_n)  //  output,  width = 1, out_reset.reset_n
	);

	qsys_top_iopll_0 ftile_iopll_ptp_sampling (
		.refclk   (ftile_iopll_ptp_sampling_refclk_clk),  //   input,  width = 1,  refclk.clk
		.locked   (),                                     //  output,  width = 1,  locked.export
		.rst      (ftile_iopll_ptp_sampling_reset_reset), //   input,  width = 1,   reset.reset
		.outclk_0 (ftile_iopll_ptp_sampling_outclk0_clk)  //  output,  width = 1, outclk0.clk
	);

	ftile_iopll_todsync_sampling ftile_iopll_todsync_sampling (
		.refclk   (ftile_iopll_todsync_sampling_refclk_clk),  //   input,  width = 1,  refclk.clk
		.locked   (ftile_iopll_todsync_sampling_locked_lock), //  output,  width = 1,  locked.lock
		.rst      (ftile_iopll_todsync_sampling_reset_reset), //   input,  width = 1,   reset.reset
		.outclk_0 (ftile_iopll_todsync_sampling_outclk0_clk)  //  output,  width = 1, outclk0.clk
	);

	qsys_top_master_todclk_0 qsys_top_master_todclk_0 (
		.in_clk  (qsys_top_master_todclk_0_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (qsys_top_master_todclk_0_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	rst_in rst_in (
		.clk         (rst_in_clk_clk),           //   input,  width = 1,       clk.clk
		.in_reset_n  (rst_in_in_reset_reset_n),  //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (rst_in_out_reset_reset_n)  //  output,  width = 1, out_reset.reset_n
	);

	sysid sysid (
		.clock    (sysid_clk_clk),                //   input,   width = 1,           clk.clk
		.reset_n  (sysid_reset_reset_n),          //   input,   width = 1,         reset.reset_n
		.readdata (sysid_control_slave_readdata), //  output,  width = 32, control_slave.readdata
		.address  (sysid_control_slave_address)   //   input,   width = 1,              .address
	);

	user_rst_clkgate_0 user_rst_clkgate_0 (
		.ninit_done (user_rst_clkgate_0_ninit_done_ninit_done)  //  output,  width = 1, ninit_done.ninit_done
	);

endmodule
