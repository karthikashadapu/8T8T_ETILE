// j204c_f_rx_tx_ip.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module j204c_f_rx_tx_ip (
		input  wire [20:0]  intel_jesd204c_f_reconfig_xcvr_address,        //         intel_jesd204c_f_reconfig_xcvr.address
		input  wire         intel_jesd204c_f_reconfig_xcvr_read,           //                                       .read
		input  wire         intel_jesd204c_f_reconfig_xcvr_write,          //                                       .write
		input  wire [31:0]  intel_jesd204c_f_reconfig_xcvr_writedata,      //                                       .writedata
		output wire [31:0]  intel_jesd204c_f_reconfig_xcvr_readdata,       //                                       .readdata
		output wire         intel_jesd204c_f_reconfig_xcvr_waitrequest,    //                                       .waitrequest
		input  wire [3:0]   intel_jesd204c_f_reconfig_xcvr_byteenable,     //                                       .byteenable
		output wire         intel_jesd204c_f_j204c_tx_rst_ack_n_export,    //    intel_jesd204c_f_j204c_tx_rst_ack_n.export
		input  wire         intel_jesd204c_f_j204c_txlclk_ctrl_export,     //     intel_jesd204c_f_j204c_txlclk_ctrl.export
		input  wire         intel_jesd204c_f_j204c_txfclk_ctrl_export,     //     intel_jesd204c_f_j204c_txfclk_ctrl.export
		input  wire         intel_jesd204c_f_j204c_tx_avs_chipselect,      //          intel_jesd204c_f_j204c_tx_avs.chipselect
		input  wire [9:0]   intel_jesd204c_f_j204c_tx_avs_address,         //                                       .address
		input  wire         intel_jesd204c_f_j204c_tx_avs_read,            //                                       .read
		output wire [31:0]  intel_jesd204c_f_j204c_tx_avs_readdata,        //                                       .readdata
		output wire         intel_jesd204c_f_j204c_tx_avs_waitrequest,     //                                       .waitrequest
		input  wire         intel_jesd204c_f_j204c_tx_avs_write,           //                                       .write
		input  wire [31:0]  intel_jesd204c_f_j204c_tx_avs_writedata,       //                                       .writedata
		input  wire [511:0] intel_jesd204c_f_j204c_tx_avst_data,           //         intel_jesd204c_f_j204c_tx_avst.data
		input  wire         intel_jesd204c_f_j204c_tx_avst_valid,          //                                       .valid
		output wire         intel_jesd204c_f_j204c_tx_avst_ready,          //                                       .ready
		input  wire         intel_jesd204c_f_j204c_tx_avst_control_export, // intel_jesd204c_f_j204c_tx_avst_control.export
		input  wire [47:0]  intel_jesd204c_f_j204c_tx_cmd_data,            //          intel_jesd204c_f_j204c_tx_cmd.data
		input  wire         intel_jesd204c_f_j204c_tx_cmd_valid,           //                                       .valid
		output wire         intel_jesd204c_f_j204c_tx_cmd_ready,           //                                       .ready
		input  wire         intel_jesd204c_f_j204c_tx_sysref_export,       //       intel_jesd204c_f_j204c_tx_sysref.export
		output wire [3:0]   intel_jesd204c_f_j204c_tx_csr_l_export,        //        intel_jesd204c_f_j204c_tx_csr_l.export
		output wire [7:0]   intel_jesd204c_f_j204c_tx_csr_f_export,        //        intel_jesd204c_f_j204c_tx_csr_f.export
		output wire [7:0]   intel_jesd204c_f_j204c_tx_csr_m_export,        //        intel_jesd204c_f_j204c_tx_csr_m.export
		output wire [1:0]   intel_jesd204c_f_j204c_tx_csr_cs_export,       //       intel_jesd204c_f_j204c_tx_csr_cs.export
		output wire [4:0]   intel_jesd204c_f_j204c_tx_csr_n_export,        //        intel_jesd204c_f_j204c_tx_csr_n.export
		output wire [4:0]   intel_jesd204c_f_j204c_tx_csr_np_export,       //       intel_jesd204c_f_j204c_tx_csr_np.export
		output wire [4:0]   intel_jesd204c_f_j204c_tx_csr_s_export,        //        intel_jesd204c_f_j204c_tx_csr_s.export
		output wire         intel_jesd204c_f_j204c_tx_csr_hd_export,       //       intel_jesd204c_f_j204c_tx_csr_hd.export
		output wire [4:0]   intel_jesd204c_f_j204c_tx_csr_cf_export,       //       intel_jesd204c_f_j204c_tx_csr_cf.export
		output wire [7:0]   intel_jesd204c_f_j204c_tx_csr_e_export,        //        intel_jesd204c_f_j204c_tx_csr_e.export
		output wire         intel_jesd204c_f_j204c_tx_int_irq,             //          intel_jesd204c_f_j204c_tx_int.irq
		input  wire         intel_jesd204c_f_j204c_rx_avs_chipselect,      //          intel_jesd204c_f_j204c_rx_avs.chipselect
		input  wire [9:0]   intel_jesd204c_f_j204c_rx_avs_address,         //                                       .address
		input  wire         intel_jesd204c_f_j204c_rx_avs_read,            //                                       .read
		output wire [31:0]  intel_jesd204c_f_j204c_rx_avs_readdata,        //                                       .readdata
		output wire         intel_jesd204c_f_j204c_rx_avs_waitrequest,     //                                       .waitrequest
		input  wire         intel_jesd204c_f_j204c_rx_avs_write,           //                                       .write
		input  wire [31:0]  intel_jesd204c_f_j204c_rx_avs_writedata,       //                                       .writedata
		output wire         intel_jesd204c_f_j204c_rx_int_irq,             //          intel_jesd204c_f_j204c_rx_int.irq
		output wire [3:0]   intel_jesd204c_f_j204c_rx_csr_l_export,        //        intel_jesd204c_f_j204c_rx_csr_l.export
		output wire [7:0]   intel_jesd204c_f_j204c_rx_csr_f_export,        //        intel_jesd204c_f_j204c_rx_csr_f.export
		output wire [7:0]   intel_jesd204c_f_j204c_rx_csr_m_export,        //        intel_jesd204c_f_j204c_rx_csr_m.export
		output wire [1:0]   intel_jesd204c_f_j204c_rx_csr_cs_export,       //       intel_jesd204c_f_j204c_rx_csr_cs.export
		output wire [4:0]   intel_jesd204c_f_j204c_rx_csr_n_export,        //        intel_jesd204c_f_j204c_rx_csr_n.export
		output wire [4:0]   intel_jesd204c_f_j204c_rx_csr_np_export,       //       intel_jesd204c_f_j204c_rx_csr_np.export
		output wire [4:0]   intel_jesd204c_f_j204c_rx_csr_s_export,        //        intel_jesd204c_f_j204c_rx_csr_s.export
		output wire         intel_jesd204c_f_j204c_rx_csr_hd_export,       //       intel_jesd204c_f_j204c_rx_csr_hd.export
		output wire [4:0]   intel_jesd204c_f_j204c_rx_csr_cf_export,       //       intel_jesd204c_f_j204c_rx_csr_cf.export
		output wire [7:0]   intel_jesd204c_f_j204c_rx_csr_e_export,        //        intel_jesd204c_f_j204c_rx_csr_e.export
		output wire [1:0]   intel_jesd204c_f_j204c_rx_csr_testmode_export, // intel_jesd204c_f_j204c_rx_csr_testmode.export
		input  wire         intel_jesd204c_f_j204c_rxlclk_ctrl_export,     //     intel_jesd204c_f_j204c_rxlclk_ctrl.export
		input  wire         intel_jesd204c_f_j204c_rxfclk_ctrl_export,     //     intel_jesd204c_f_j204c_rxfclk_ctrl.export
		input  wire         intel_jesd204c_f_j204c_rx_sysref_export,       //       intel_jesd204c_f_j204c_rx_sysref.export
		output wire         intel_jesd204c_f_j204c_rx_rst_ack_n_export,    //    intel_jesd204c_f_j204c_rx_rst_ack_n.export
		output wire [511:0] intel_jesd204c_f_j204c_rx_avst_data,           //         intel_jesd204c_f_j204c_rx_avst.data
		output wire         intel_jesd204c_f_j204c_rx_avst_valid,          //                                       .valid
		input  wire         intel_jesd204c_f_j204c_rx_avst_ready,          //                                       .ready
		output wire         intel_jesd204c_f_j204c_rx_avst_control_export, // intel_jesd204c_f_j204c_rx_avst_control.export
		output wire [47:0]  intel_jesd204c_f_j204c_rx_cmd_data,            //          intel_jesd204c_f_j204c_rx_cmd.data
		output wire         intel_jesd204c_f_j204c_rx_cmd_valid,           //                                       .valid
		input  wire         intel_jesd204c_f_j204c_rx_cmd_ready,           //                                       .ready
		output wire [7:0]   intel_jesd204c_f_j204c_rx_cmd_par_err_export,  //  intel_jesd204c_f_j204c_rx_cmd_par_err.export
		output wire         intel_jesd204c_f_j204c_rx_sh_lock_export,      //      intel_jesd204c_f_j204c_rx_sh_lock.export
		output wire         intel_jesd204c_f_j204c_rx_emb_lock_export,     //     intel_jesd204c_f_j204c_rx_emb_lock.export
		output wire [7:0]   intel_jesd204c_f_j204c_rx_crc_err_export,      //      intel_jesd204c_f_j204c_rx_crc_err.export
		output wire [7:0]   intel_jesd204c_f_tx_serial_data_export,        //        intel_jesd204c_f_tx_serial_data.export
		output wire [7:0]   intel_jesd204c_f_tx_serial_data_n_export,      //      intel_jesd204c_f_tx_serial_data_n.export
		input  wire [7:0]   intel_jesd204c_f_rx_serial_data_export,        //        intel_jesd204c_f_rx_serial_data.export
		input  wire [7:0]   intel_jesd204c_f_rx_serial_data_n_export,      //      intel_jesd204c_f_rx_serial_data_n.export
		input  wire         jesd_link_clk_in_clk_clk,                      //                   jesd_link_clk_in_clk.clk
		input  wire         mgmt_clk_in_clk_clk,                           //                        mgmt_clk_in_clk.clk
		input  wire         mgmt_reset_in_reset_reset_n,                   //                    mgmt_reset_in_reset.reset_n
		output wire         reset_out1_reset,                              //                             reset_out1.reset
		output wire         reset_out2_reset,                              //                             reset_out2.reset
		output wire         reset_out4_reset,                              //                             reset_out4.reset
		input  wire         reset1_dsrt_qual_reset1_dsrt_qual,             //                       reset1_dsrt_qual.reset1_dsrt_qual
		input  wire         reset2_dsrt_qual_reset2_dsrt_qual,             //                       reset2_dsrt_qual.reset2_dsrt_qual
		input  wire         reset4_dsrt_qual_reset4_dsrt_qual,             //                       reset4_dsrt_qual.reset4_dsrt_qual
		input  wire [7:0]   reset_sequencer_0_av_csr_address,              //               reset_sequencer_0_av_csr.address
		output wire [31:0]  reset_sequencer_0_av_csr_readdata,             //                                       .readdata
		input  wire         reset_sequencer_0_av_csr_read,                 //                                       .read
		input  wire [31:0]  reset_sequencer_0_av_csr_writedata,            //                                       .writedata
		input  wire         reset_sequencer_0_av_csr_write,                //                                       .write
		output wire         reset_sequencer_0_av_csr_irq_irq,              //           reset_sequencer_0_av_csr_irq.irq
		input  wire         systemclk_f_refclk_fgt_in_refclk_fgt_0         //                 systemclk_f_refclk_fgt.in_refclk_fgt_0
	);

	wire    mgmt_clk_out_clk_clk;                            // mgmt_clk:out_clk -> [avs_reset:clk, intel_jesd204c_f:j204c_rx_avs_clk, intel_jesd204c_f:j204c_tx_avs_clk, intel_jesd204c_f:reconfig_xcvr_clk, mgmt_reset:clk, reset_controller_0:clk, reset_sequencer_0:clk, rx_reset:clk, tx_reset:clk]
	wire    jesd_link_clk_out_clk_clk;                       // jesd_link_clk:out_clk -> [intel_jesd204c_f:j204c_rxframe_clk, intel_jesd204c_f:j204c_rxlink_clk, intel_jesd204c_f:j204c_txframe_clk, intel_jesd204c_f:j204c_txlink_clk]
	wire    intel_jesd204c_f_j204c_rx_dev_lane_align_export; // intel_jesd204c_f:j204c_rx_dev_lane_align -> intel_jesd204c_f:j204c_rx_alldev_lane_align
	wire    systemclk_f_out_refclk_fgt_0_clk;                // systemclk_f:out_refclk_fgt_0 -> intel_jesd204c_f:j204c_pll_refclk
	wire    systemclk_f_out_systempll_clk_0_clk;             // systemclk_f:out_systempll_clk_0 -> intel_jesd204c_f:sysclk
	wire    mgmt_reset_out_reset_reset;                      // mgmt_reset:out_reset_n -> [intel_jesd204c_f:reconfig_xcvr_reset, reset_controller_0:reset_in0, reset_sequencer_0:csr_reset, reset_sequencer_0:reset_in0]
	wire    avs_reset_out_reset_reset;                       // avs_reset:out_reset_n -> [intel_jesd204c_f:j204c_rx_avs_rst_n, intel_jesd204c_f:j204c_tx_avs_rst_n]
	wire    rx_reset_out_reset_reset;                        // rx_reset:out_reset_n -> intel_jesd204c_f:j204c_rx_rst_n
	wire    tx_reset_out_reset_reset;                        // tx_reset:out_reset_n -> intel_jesd204c_f:j204c_tx_rst_n
	wire    reset_sequencer_0_reset_out0_reset;              // reset_sequencer_0:reset_out0 -> avs_reset:in_reset_n
	wire    reset_sequencer_0_reset_out3_reset;              // reset_sequencer_0:reset_out3 -> tx_reset:in_reset_n
	wire    reset_sequencer_0_reset_out5_reset;              // reset_sequencer_0:reset_out5 -> rx_reset:in_reset_n

	j204c_f_rx_tx_ip_reset_bridge_2 avs_reset (
		.clk         (mgmt_clk_out_clk_clk),                //   input,  width = 1,       clk.clk
		.in_reset_n  (~reset_sequencer_0_reset_out0_reset), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (avs_reset_out_reset_reset)            //  output,  width = 1, out_reset.reset_n
	);

	j204c_f_rx_tx_ip_intel_jesd204c_f intel_jesd204c_f (
		.reconfig_xcvr_clk          (mgmt_clk_out_clk_clk),                            //   input,    width = 1,          reconfig_xcvr_clk.clk
		.reconfig_xcvr_reset        (~mgmt_reset_out_reset_reset),                     //   input,    width = 1,        reconfig_xcvr_reset.reset
		.reconfig_xcvr_address      (intel_jesd204c_f_reconfig_xcvr_address),          //   input,   width = 21,              reconfig_xcvr.address
		.reconfig_xcvr_read         (intel_jesd204c_f_reconfig_xcvr_read),             //   input,    width = 1,                           .read
		.reconfig_xcvr_write        (intel_jesd204c_f_reconfig_xcvr_write),            //   input,    width = 1,                           .write
		.reconfig_xcvr_writedata    (intel_jesd204c_f_reconfig_xcvr_writedata),        //   input,   width = 32,                           .writedata
		.reconfig_xcvr_readdata     (intel_jesd204c_f_reconfig_xcvr_readdata),         //  output,   width = 32,                           .readdata
		.reconfig_xcvr_waitrequest  (intel_jesd204c_f_reconfig_xcvr_waitrequest),      //  output,    width = 1,                           .waitrequest
		.reconfig_xcvr_byteenable   (intel_jesd204c_f_reconfig_xcvr_byteenable),       //   input,    width = 4,                           .byteenable
		.j204c_txlink_clk           (jesd_link_clk_out_clk_clk),                       //   input,    width = 1,           j204c_txlink_clk.clk
		.j204c_txframe_clk          (jesd_link_clk_out_clk_clk),                       //   input,    width = 1,          j204c_txframe_clk.clk
		.j204c_tx_rst_n             (tx_reset_out_reset_reset),                        //   input,    width = 1,             j204c_tx_rst_n.reset_n
		.j204c_tx_rst_ack_n         (intel_jesd204c_f_j204c_tx_rst_ack_n_export),      //  output,    width = 1,         j204c_tx_rst_ack_n.export
		.j204c_txlclk_ctrl          (intel_jesd204c_f_j204c_txlclk_ctrl_export),       //   input,    width = 1,          j204c_txlclk_ctrl.export
		.j204c_txfclk_ctrl          (intel_jesd204c_f_j204c_txfclk_ctrl_export),       //   input,    width = 1,          j204c_txfclk_ctrl.export
		.j204c_tx_avs_clk           (mgmt_clk_out_clk_clk),                            //   input,    width = 1,           j204c_tx_avs_clk.clk
		.j204c_tx_avs_rst_n         (avs_reset_out_reset_reset),                       //   input,    width = 1,         j204c_tx_avs_rst_n.reset_n
		.j204c_tx_avs_chipselect    (intel_jesd204c_f_j204c_tx_avs_chipselect),        //   input,    width = 1,               j204c_tx_avs.chipselect
		.j204c_tx_avs_address       (intel_jesd204c_f_j204c_tx_avs_address),           //   input,   width = 10,                           .address
		.j204c_tx_avs_read          (intel_jesd204c_f_j204c_tx_avs_read),              //   input,    width = 1,                           .read
		.j204c_tx_avs_readdata      (intel_jesd204c_f_j204c_tx_avs_readdata),          //  output,   width = 32,                           .readdata
		.j204c_tx_avs_waitrequest   (intel_jesd204c_f_j204c_tx_avs_waitrequest),       //  output,    width = 1,                           .waitrequest
		.j204c_tx_avs_write         (intel_jesd204c_f_j204c_tx_avs_write),             //   input,    width = 1,                           .write
		.j204c_tx_avs_writedata     (intel_jesd204c_f_j204c_tx_avs_writedata),         //   input,   width = 32,                           .writedata
		.j204c_tx_avst_data         (intel_jesd204c_f_j204c_tx_avst_data),             //   input,  width = 512,              j204c_tx_avst.data
		.j204c_tx_avst_valid        (intel_jesd204c_f_j204c_tx_avst_valid),            //   input,    width = 1,                           .valid
		.j204c_tx_avst_ready        (intel_jesd204c_f_j204c_tx_avst_ready),            //  output,    width = 1,                           .ready
		.j204c_tx_avst_control      (intel_jesd204c_f_j204c_tx_avst_control_export),   //   input,    width = 1,      j204c_tx_avst_control.export
		.j204c_tx_cmd_data          (intel_jesd204c_f_j204c_tx_cmd_data),              //   input,   width = 48,               j204c_tx_cmd.data
		.j204c_tx_cmd_valid         (intel_jesd204c_f_j204c_tx_cmd_valid),             //   input,    width = 1,                           .valid
		.j204c_tx_cmd_ready         (intel_jesd204c_f_j204c_tx_cmd_ready),             //  output,    width = 1,                           .ready
		.j204c_tx_sysref            (intel_jesd204c_f_j204c_tx_sysref_export),         //   input,    width = 1,            j204c_tx_sysref.export
		.j204c_tx_csr_l             (intel_jesd204c_f_j204c_tx_csr_l_export),          //  output,    width = 4,             j204c_tx_csr_l.export
		.j204c_tx_csr_f             (intel_jesd204c_f_j204c_tx_csr_f_export),          //  output,    width = 8,             j204c_tx_csr_f.export
		.j204c_tx_csr_m             (intel_jesd204c_f_j204c_tx_csr_m_export),          //  output,    width = 8,             j204c_tx_csr_m.export
		.j204c_tx_csr_cs            (intel_jesd204c_f_j204c_tx_csr_cs_export),         //  output,    width = 2,            j204c_tx_csr_cs.export
		.j204c_tx_csr_n             (intel_jesd204c_f_j204c_tx_csr_n_export),          //  output,    width = 5,             j204c_tx_csr_n.export
		.j204c_tx_csr_np            (intel_jesd204c_f_j204c_tx_csr_np_export),         //  output,    width = 5,            j204c_tx_csr_np.export
		.j204c_tx_csr_s             (intel_jesd204c_f_j204c_tx_csr_s_export),          //  output,    width = 5,             j204c_tx_csr_s.export
		.j204c_tx_csr_hd            (intel_jesd204c_f_j204c_tx_csr_hd_export),         //  output,    width = 1,            j204c_tx_csr_hd.export
		.j204c_tx_csr_cf            (intel_jesd204c_f_j204c_tx_csr_cf_export),         //  output,    width = 5,            j204c_tx_csr_cf.export
		.j204c_tx_csr_e             (intel_jesd204c_f_j204c_tx_csr_e_export),          //  output,    width = 8,             j204c_tx_csr_e.export
		.j204c_tx_int               (intel_jesd204c_f_j204c_tx_int_irq),               //  output,    width = 1,               j204c_tx_int.irq
		.j204c_rx_avs_clk           (mgmt_clk_out_clk_clk),                            //   input,    width = 1,           j204c_rx_avs_clk.clk
		.j204c_rx_avs_rst_n         (avs_reset_out_reset_reset),                       //   input,    width = 1,         j204c_rx_avs_rst_n.reset_n
		.j204c_rx_avs_chipselect    (intel_jesd204c_f_j204c_rx_avs_chipselect),        //   input,    width = 1,               j204c_rx_avs.chipselect
		.j204c_rx_avs_address       (intel_jesd204c_f_j204c_rx_avs_address),           //   input,   width = 10,                           .address
		.j204c_rx_avs_read          (intel_jesd204c_f_j204c_rx_avs_read),              //   input,    width = 1,                           .read
		.j204c_rx_avs_readdata      (intel_jesd204c_f_j204c_rx_avs_readdata),          //  output,   width = 32,                           .readdata
		.j204c_rx_avs_waitrequest   (intel_jesd204c_f_j204c_rx_avs_waitrequest),       //  output,    width = 1,                           .waitrequest
		.j204c_rx_avs_write         (intel_jesd204c_f_j204c_rx_avs_write),             //   input,    width = 1,                           .write
		.j204c_rx_avs_writedata     (intel_jesd204c_f_j204c_rx_avs_writedata),         //   input,   width = 32,                           .writedata
		.j204c_rx_int               (intel_jesd204c_f_j204c_rx_int_irq),               //  output,    width = 1,               j204c_rx_int.irq
		.j204c_rx_csr_l             (intel_jesd204c_f_j204c_rx_csr_l_export),          //  output,    width = 4,             j204c_rx_csr_l.export
		.j204c_rx_csr_f             (intel_jesd204c_f_j204c_rx_csr_f_export),          //  output,    width = 8,             j204c_rx_csr_f.export
		.j204c_rx_csr_m             (intel_jesd204c_f_j204c_rx_csr_m_export),          //  output,    width = 8,             j204c_rx_csr_m.export
		.j204c_rx_csr_cs            (intel_jesd204c_f_j204c_rx_csr_cs_export),         //  output,    width = 2,            j204c_rx_csr_cs.export
		.j204c_rx_csr_n             (intel_jesd204c_f_j204c_rx_csr_n_export),          //  output,    width = 5,             j204c_rx_csr_n.export
		.j204c_rx_csr_np            (intel_jesd204c_f_j204c_rx_csr_np_export),         //  output,    width = 5,            j204c_rx_csr_np.export
		.j204c_rx_csr_s             (intel_jesd204c_f_j204c_rx_csr_s_export),          //  output,    width = 5,             j204c_rx_csr_s.export
		.j204c_rx_csr_hd            (intel_jesd204c_f_j204c_rx_csr_hd_export),         //  output,    width = 1,            j204c_rx_csr_hd.export
		.j204c_rx_csr_cf            (intel_jesd204c_f_j204c_rx_csr_cf_export),         //  output,    width = 5,            j204c_rx_csr_cf.export
		.j204c_rx_csr_e             (intel_jesd204c_f_j204c_rx_csr_e_export),          //  output,    width = 8,             j204c_rx_csr_e.export
		.j204c_rx_csr_testmode      (intel_jesd204c_f_j204c_rx_csr_testmode_export),   //  output,    width = 2,      j204c_rx_csr_testmode.export
		.j204c_rxlink_clk           (jesd_link_clk_out_clk_clk),                       //   input,    width = 1,           j204c_rxlink_clk.clk
		.j204c_rxframe_clk          (jesd_link_clk_out_clk_clk),                       //   input,    width = 1,          j204c_rxframe_clk.clk
		.j204c_rxlclk_ctrl          (intel_jesd204c_f_j204c_rxlclk_ctrl_export),       //   input,    width = 1,          j204c_rxlclk_ctrl.export
		.j204c_rxfclk_ctrl          (intel_jesd204c_f_j204c_rxfclk_ctrl_export),       //   input,    width = 1,          j204c_rxfclk_ctrl.export
		.j204c_rx_sysref            (intel_jesd204c_f_j204c_rx_sysref_export),         //   input,    width = 1,            j204c_rx_sysref.export
		.j204c_rx_rst_n             (rx_reset_out_reset_reset),                        //   input,    width = 1,             j204c_rx_rst_n.reset_n
		.j204c_rx_rst_ack_n         (intel_jesd204c_f_j204c_rx_rst_ack_n_export),      //  output,    width = 1,         j204c_rx_rst_ack_n.export
		.j204c_rx_alldev_lane_align (intel_jesd204c_f_j204c_rx_dev_lane_align_export), //   input,    width = 1, j204c_rx_alldev_lane_align.export
		.j204c_rx_dev_lane_align    (intel_jesd204c_f_j204c_rx_dev_lane_align_export), //  output,    width = 1,    j204c_rx_dev_lane_align.export
		.j204c_rx_avst_data         (intel_jesd204c_f_j204c_rx_avst_data),             //  output,  width = 512,              j204c_rx_avst.data
		.j204c_rx_avst_valid        (intel_jesd204c_f_j204c_rx_avst_valid),            //  output,    width = 1,                           .valid
		.j204c_rx_avst_ready        (intel_jesd204c_f_j204c_rx_avst_ready),            //   input,    width = 1,                           .ready
		.j204c_rx_avst_control      (intel_jesd204c_f_j204c_rx_avst_control_export),   //  output,    width = 1,      j204c_rx_avst_control.export
		.j204c_rx_cmd_data          (intel_jesd204c_f_j204c_rx_cmd_data),              //  output,   width = 48,               j204c_rx_cmd.data
		.j204c_rx_cmd_valid         (intel_jesd204c_f_j204c_rx_cmd_valid),             //  output,    width = 1,                           .valid
		.j204c_rx_cmd_ready         (intel_jesd204c_f_j204c_rx_cmd_ready),             //   input,    width = 1,                           .ready
		.j204c_rx_cmd_par_err       (intel_jesd204c_f_j204c_rx_cmd_par_err_export),    //  output,    width = 8,       j204c_rx_cmd_par_err.export
		.j204c_rx_sh_lock           (intel_jesd204c_f_j204c_rx_sh_lock_export),        //  output,    width = 1,           j204c_rx_sh_lock.export
		.j204c_rx_emb_lock          (intel_jesd204c_f_j204c_rx_emb_lock_export),       //  output,    width = 1,          j204c_rx_emb_lock.export
		.j204c_rx_crc_err           (intel_jesd204c_f_j204c_rx_crc_err_export),        //  output,    width = 8,           j204c_rx_crc_err.export
		.j204c_syspll_div2_clk      (),                                                //  output,    width = 1,      j204c_syspll_div2_clk.export
		.j204c_pll_refclk           (systemclk_f_out_refclk_fgt_0_clk),                //   input,    width = 1,           j204c_pll_refclk.clk
		.sysclk                     (systemclk_f_out_systempll_clk_0_clk),             //   input,    width = 1,                     sysclk.clk
		.tx_serial_data             (intel_jesd204c_f_tx_serial_data_export),          //  output,    width = 8,             tx_serial_data.export
		.tx_serial_data_n           (intel_jesd204c_f_tx_serial_data_n_export),        //  output,    width = 8,           tx_serial_data_n.export
		.rx_serial_data             (intel_jesd204c_f_rx_serial_data_export),          //   input,    width = 8,             rx_serial_data.export
		.rx_serial_data_n           (intel_jesd204c_f_rx_serial_data_n_export)         //   input,    width = 8,           rx_serial_data_n.export
	);

	j204c_f_rx_tx_ip_clock_bridge_1 jesd_link_clk (
		.in_clk  (jesd_link_clk_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (jesd_link_clk_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	j204c_f_rx_tx_ip_clock_bridge_0 mgmt_clk (
		.in_clk  (mgmt_clk_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (mgmt_clk_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	j204c_f_rx_tx_ip_reset_bridge_0 mgmt_reset (
		.clk         (mgmt_clk_out_clk_clk),        //   input,  width = 1,       clk.clk
		.in_reset_n  (mgmt_reset_in_reset_reset_n), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (mgmt_reset_out_reset_reset)   //  output,  width = 1, out_reset.reset_n
	);

	j204c_f_rx_tx_ip_reset_controller_0 reset_controller_0 (
		.reset_in0 (~mgmt_reset_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk       (mgmt_clk_out_clk_clk),        //   input,  width = 1,       clk.clk
		.reset_out ()                             //  output,  width = 1, reset_out.reset
	);

	j204c_f_rx_tx_ip_reset_sequencer_0 reset_sequencer_0 (
		.clk              (mgmt_clk_out_clk_clk),               //   input,   width = 1,              clk.clk
		.reset_in0        (~mgmt_reset_out_reset_reset),        //   input,   width = 1,        reset_in0.reset
		.reset_out0       (reset_sequencer_0_reset_out0_reset), //  output,   width = 1,       reset_out0.reset
		.reset_out1       (reset_out1_reset),                   //  output,   width = 1,       reset_out1.reset
		.reset_out2       (reset_out2_reset),                   //  output,   width = 1,       reset_out2.reset
		.reset_out3       (reset_sequencer_0_reset_out3_reset), //  output,   width = 1,       reset_out3.reset
		.reset_out4       (reset_out4_reset),                   //  output,   width = 1,       reset_out4.reset
		.reset_out5       (reset_sequencer_0_reset_out5_reset), //  output,   width = 1,       reset_out5.reset
		.reset1_dsrt_qual (reset1_dsrt_qual_reset1_dsrt_qual),  //   input,   width = 1, reset1_dsrt_qual.reset1_dsrt_qual
		.reset2_dsrt_qual (reset2_dsrt_qual_reset2_dsrt_qual),  //   input,   width = 1, reset2_dsrt_qual.reset2_dsrt_qual
		.reset4_dsrt_qual (reset4_dsrt_qual_reset4_dsrt_qual),  //   input,   width = 1, reset4_dsrt_qual.reset4_dsrt_qual
		.csr_reset        (~mgmt_reset_out_reset_reset),        //   input,   width = 1,        csr_reset.reset
		.av_address       (reset_sequencer_0_av_csr_address),   //   input,   width = 8,           av_csr.address
		.av_readdata      (reset_sequencer_0_av_csr_readdata),  //  output,  width = 32,                 .readdata
		.av_read          (reset_sequencer_0_av_csr_read),      //   input,   width = 1,                 .read
		.av_writedata     (reset_sequencer_0_av_csr_writedata), //   input,  width = 32,                 .writedata
		.av_write         (reset_sequencer_0_av_csr_write),     //   input,   width = 1,                 .write
		.irq              (reset_sequencer_0_av_csr_irq_irq)    //  output,   width = 1,       av_csr_irq.irq
	);

	j204c_f_rx_tx_ip_tx_reset_0 rx_reset (
		.clk         (mgmt_clk_out_clk_clk),                //   input,  width = 1,       clk.clk
		.in_reset_n  (~reset_sequencer_0_reset_out5_reset), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (rx_reset_out_reset_reset)             //  output,  width = 1, out_reset.reset_n
	);

	j204c_f_rx_tx_ip_systemclk_f systemclk_f (
		.out_systempll_synthlock_0 (),                                       //  output,  width = 1, out_systempll_synthlock_0.out_systempll_synthlock
		.out_systempll_clk_0       (systemclk_f_out_systempll_clk_0_clk),    //  output,  width = 1,       out_systempll_clk_0.clk
		.out_refclk_fgt_0          (systemclk_f_out_refclk_fgt_0_clk),       //  output,  width = 1,          out_refclk_fgt_0.clk
		.in_refclk_fgt_0           (systemclk_f_refclk_fgt_in_refclk_fgt_0)  //   input,  width = 1,                refclk_fgt.in_refclk_fgt_0
	);

	j204c_f_rx_tx_ip_avs_reset_0 tx_reset (
		.clk         (mgmt_clk_out_clk_clk),                //   input,  width = 1,       clk.clk
		.in_reset_n  (~reset_sequencer_0_reset_out3_reset), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (tx_reset_out_reset_reset)             //  output,  width = 1, out_reset.reset_n
	);

endmodule
