// master_tod_subsys.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module master_tod_subsys (
		input  wire        master_tod_top_0_csr_write,                                //                       master_tod_top_0_csr.write
		input  wire [31:0] master_tod_top_0_csr_writedata,                            //                                           .writedata
		input  wire        master_tod_top_0_csr_read,                                 //                                           .read
		output wire [31:0] master_tod_top_0_csr_readdata,                             //                                           .readdata
		output wire        master_tod_top_0_csr_waitrequest,                          //                                           .waitrequest
		input  wire [3:0]  master_tod_top_0_csr_address,                              //                                           .address
		input  wire        master_tod_top_0_i_clk_tod_clk,                            //                 master_tod_top_0_i_clk_tod.clk
		input  wire        master_tod_top_0_i_reconfig_rst_n_reset_n,                 //          master_tod_top_0_i_reconfig_rst_n.reset_n
		input  wire        master_tod_top_0_i_tod_rst_n_reset_n,                      //               master_tod_top_0_i_tod_rst_n.reset_n
		output wire        master_tod_top_0_pulse_per_second_pps,                     //          master_tod_top_0_pulse_per_second.pps
		output wire        master_tod_top_0_avst_tod_data_valid,                      //             master_tod_top_0_avst_tod_data.valid
		output wire [95:0] master_tod_top_0_avst_tod_data_data,                       //                                           .data
		input  wire        master_tod_top_0_i_upstr_pll_lock,                         //               master_tod_top_0_i_upstr_pll.lock
		input  wire        mtod_subsys_clk100_in_clk_clk,                             //                  mtod_subsys_clk100_in_clk.clk
		input  wire        mtod_subsys_pps_load_tod_0_period_clock_clk,               //    mtod_subsys_pps_load_tod_0_period_clock.clk
		input  wire        mtod_subsys_pps_load_tod_0_reset_reset,                    //           mtod_subsys_pps_load_tod_0_reset.reset
		input  wire        mtod_subsys_pps_load_tod_0_csr_reset_reset,                //       mtod_subsys_pps_load_tod_0_csr_reset.reset
		output wire [31:0] mtod_subsys_pps_load_tod_0_csr_readdata,                   //             mtod_subsys_pps_load_tod_0_csr.readdata
		input  wire        mtod_subsys_pps_load_tod_0_csr_write,                      //                                           .write
		input  wire        mtod_subsys_pps_load_tod_0_csr_read,                       //                                           .read
		input  wire [31:0] mtod_subsys_pps_load_tod_0_csr_writedata,                  //                                           .writedata
		output wire        mtod_subsys_pps_load_tod_0_csr_waitrequest,                //                                           .waitrequest
		input  wire [5:0]  mtod_subsys_pps_load_tod_0_csr_address,                    //                                           .address
		input  wire        mtod_subsys_pps_load_tod_0_pps_interface_pulse_per_second, //   mtod_subsys_pps_load_tod_0_pps_interface.pulse_per_second
		input  wire [95:0] mtod_subsys_pps_load_tod_0_time_of_day_96b_data,           // mtod_subsys_pps_load_tod_0_time_of_day_96b.data
		output wire        mtod_subsys_pps_load_tod_0_pps_irq_irq,                    //         mtod_subsys_pps_load_tod_0_pps_irq.irq
		input  wire        mtod_subsys_rstn_in_reset_reset_n                          //                  mtod_subsys_rstn_in_reset.reset_n
	);

	wire         mtod_subsys_clk100_out_clk_clk;                         // mtod_subsys_clk100:out_clk -> [master_tod_top_0:i_clk_reconfig, mtod_subsys_pps_load_tod_0:csr_clock, mtod_subsys_rstn:clk]
	wire         mtod_subsys_pps_load_tod_0_time_of_data_96b_load_valid; // mtod_subsys_pps_load_tod_0:time_of_data_96b_load_valid -> master_tod_top_0:i_tod_96b_load_valid
	wire  [95:0] mtod_subsys_pps_load_tod_0_time_of_data_96b_load_data;  // mtod_subsys_pps_load_tod_0:time_of_data_96b_load_data -> master_tod_top_0:i_tod_96b_load_data

	master_tod_top_0 master_tod_top_0 (
		.i_csr_write          (master_tod_top_0_csr_write),                             //   input,   width = 1,                csr.write
		.i_csr_writedata      (master_tod_top_0_csr_writedata),                         //   input,  width = 32,                   .writedata
		.i_csr_read           (master_tod_top_0_csr_read),                              //   input,   width = 1,                   .read
		.o_csr_readdata       (master_tod_top_0_csr_readdata),                          //  output,  width = 32,                   .readdata
		.o_csr_waitrequest    (master_tod_top_0_csr_waitrequest),                       //  output,   width = 1,                   .waitrequest
		.i_csr_addr           (master_tod_top_0_csr_address),                           //   input,   width = 4,                   .address
		.i_clk_reconfig       (mtod_subsys_clk100_out_clk_clk),                         //   input,   width = 1,     i_clk_reconfig.clk
		.i_clk_tod            (master_tod_top_0_i_clk_tod_clk),                         //   input,   width = 1,          i_clk_tod.clk
		.i_reconfig_rst_n     (master_tod_top_0_i_reconfig_rst_n_reset_n),              //   input,   width = 1,   i_reconfig_rst_n.reset_n
		.i_tod_rst_n          (master_tod_top_0_i_tod_rst_n_reset_n),                   //   input,   width = 1,        i_tod_rst_n.reset_n
		.i_tod_96b_load_valid (mtod_subsys_pps_load_tod_0_time_of_data_96b_load_valid), //   input,   width = 1, avst_tod_load_data.valid
		.i_tod_96b_load_data  (mtod_subsys_pps_load_tod_0_time_of_data_96b_load_data),  //   input,  width = 96,                   .data
		.o_pps                (master_tod_top_0_pulse_per_second_pps),                  //  output,   width = 1,   pulse_per_second.pps
		.o_tod_96b_valid      (master_tod_top_0_avst_tod_data_valid),                   //  output,   width = 1,      avst_tod_data.valid
		.o_tod_96b_data       (master_tod_top_0_avst_tod_data_data),                    //  output,  width = 96,                   .data
		.i_upstr_pll_lock     (master_tod_top_0_i_upstr_pll_lock)                       //   input,   width = 1,        i_upstr_pll.lock
	);

	mtod_subsys_clk100 mtod_subsys_clk100 (
		.in_clk  (mtod_subsys_clk100_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (mtod_subsys_clk100_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	mtod_subsys_pps_load_tod_0 mtod_subsys_pps_load_tod_0 (
		.period_clock                (mtod_subsys_pps_load_tod_0_period_clock_clk),               //   input,   width = 1,          period_clock.clk
		.reset                       (mtod_subsys_pps_load_tod_0_reset_reset),                    //   input,   width = 1,                 reset.reset
		.csr_clock                   (mtod_subsys_clk100_out_clk_clk),                            //   input,   width = 1,             csr_clock.clk
		.csr_reset                   (mtod_subsys_pps_load_tod_0_csr_reset_reset),                //   input,   width = 1,             csr_reset.reset
		.csr_readdata                (mtod_subsys_pps_load_tod_0_csr_readdata),                   //  output,  width = 32,                   csr.readdata
		.csr_write                   (mtod_subsys_pps_load_tod_0_csr_write),                      //   input,   width = 1,                      .write
		.csr_read                    (mtod_subsys_pps_load_tod_0_csr_read),                       //   input,   width = 1,                      .read
		.csr_writedata               (mtod_subsys_pps_load_tod_0_csr_writedata),                  //   input,  width = 32,                      .writedata
		.csr_waitrequest             (mtod_subsys_pps_load_tod_0_csr_waitrequest),                //  output,   width = 1,                      .waitrequest
		.csr_address                 (mtod_subsys_pps_load_tod_0_csr_address),                    //   input,   width = 6,                      .address
		.pps_pulse_per_second        (mtod_subsys_pps_load_tod_0_pps_interface_pulse_per_second), //   input,   width = 1,         pps_interface.pulse_per_second
		.time_of_day_96b             (mtod_subsys_pps_load_tod_0_time_of_day_96b_data),           //   input,  width = 96,       time_of_day_96b.data
		.time_of_data_96b_load_data  (mtod_subsys_pps_load_tod_0_time_of_data_96b_load_data),     //  output,  width = 96, time_of_data_96b_load.data
		.time_of_data_96b_load_valid (mtod_subsys_pps_load_tod_0_time_of_data_96b_load_valid),    //  output,   width = 1,                      .valid
		.pps_irq                     (mtod_subsys_pps_load_tod_0_pps_irq_irq)                     //  output,   width = 1,               pps_irq.irq
	);

	mtod_subsys_rstn mtod_subsys_rstn (
		.clk         (mtod_subsys_clk100_out_clk_clk),    //   input,  width = 1,       clk.clk
		.in_reset_n  (mtod_subsys_rstn_in_reset_reset_n), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n ()                                   //  output,  width = 1, out_reset.reset_n
	);

endmodule
