// tod_slave_sub_system.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module tod_slave_sub_system (
		input  wire [95:0] master_tod_split_conduit_end_data,             //             master_tod_split_conduit_end.data
		input  wire        master_tod_split_conduit_end_valid,            //                                         .valid
		output wire [95:0] master_tod_split_conduit_end_10_data,          //          master_tod_split_conduit_end_10.data
		output wire        master_tod_split_conduit_end_10_valid,         //                                         .valid
		input  wire        oran_tod_stack_tx_clk_clk,                     //                    oran_tod_stack_tx_clk.clk
		input  wire        oran_tod_stack_rx_clk_clk,                     //                    oran_tod_stack_rx_clk.clk
		input  wire        oran_tod_stack_todsync_sample_clk_clk,         //        oran_tod_stack_todsync_sample_clk.clk
		output wire [95:0] oran_tod_stack_tx_tod_interface_tdata,         //          oran_tod_stack_tx_tod_interface.tdata
		output wire        oran_tod_stack_tx_tod_interface_tvalid,        //                                         .tvalid
		output wire [95:0] oran_tod_stack_rx_tod_interface_tdata,         //          oran_tod_stack_rx_tod_interface.tdata
		output wire        oran_tod_stack_rx_tod_interface_tvalid,        //                                         .tvalid
		input  wire        oran_tod_stack_tx_pll_locked_lock,             //             oran_tod_stack_tx_pll_locked.lock
		input  wire        port_8_tod_stack_tx_clk_clk,                   //                  port_8_tod_stack_tx_clk.clk
		input  wire        port_8_tod_stack_rx_clk_clk,                   //                  port_8_tod_stack_rx_clk.clk
		input  wire        port_8_tod_stack_todsync_sample_clk_clk,       //      port_8_tod_stack_todsync_sample_clk.clk
		output wire [95:0] port_8_tod_stack_tx_tod_interface_tdata,       //        port_8_tod_stack_tx_tod_interface.tdata
		output wire        port_8_tod_stack_tx_tod_interface_tvalid,      //                                         .tvalid
		output wire [95:0] port_8_tod_stack_rx_tod_interface_tdata,       //        port_8_tod_stack_rx_tod_interface.tdata
		output wire        port_8_tod_stack_rx_tod_interface_tvalid,      //                                         .tvalid
		input  wire        port_8_tod_stack_tx_pll_locked_lock,           //           port_8_tod_stack_tx_pll_locked.lock
		input  wire        tod_subsys_clk_100_in_clk_clk,                 //                tod_subsys_clk_100_in_clk.clk
		input  wire        tod_subsys_mtod_clk_in_clk_clk,                //               tod_subsys_mtod_clk_in_clk.clk
		input  wire        tod_subsys_rst_100_in_reset_reset_n,           //              tod_subsys_rst_100_in_reset.reset_n
		input  wire [0:0]  todsync_sample_plllock_split_conduit_end_lock  // todsync_sample_plllock_split_conduit_end.lock
	);

	wire         tod_subsys_clk_100_out_clk_clk;                  // tod_subsys_clk_100:out_clk -> [oran_tod_stack:i_reconfig_clk, port_8_tod_stack:i_reconfig_clk, tod_subsys_rst_100:clk]
	wire         tod_subsys_mtod_clk_out_clk_clk;                 // tod_subsys_mtod_clk:out_clk -> [oran_ptp2gps_conv_0:clk_tod, oran_tod_stack:i_clk_master_tod, port_8_tod_stack:i_clk_master_tod, rst_controller:clk, tod_156_reset_controller_0:clk]
	wire         master_tod_split_conduit_end_1_valid;            // master_tod_split:valid_conduit_out_1 -> port_8_tod_stack:i_ptp_master_tod_valid
	wire  [95:0] master_tod_split_conduit_end_1_data;             // master_tod_split:data_conduit_out_1 -> port_8_tod_stack:i_ptp_master_tod
	wire   [0:0] todsync_sample_plllock_split_conduit_end_1_lock; // todsync_sample_plllock_split:conduit_out_1 -> port_8_tod_stack:i_clk_todsync_sample_locked
	wire   [0:0] todsync_sample_plllock_split_conduit_end_3_lock; // todsync_sample_plllock_split:conduit_out_3 -> oran_tod_stack:i_clk_todsync_sample_locked
	wire         oran_ptp2gps_conv_0_gps_seconds_valid;           // oran_ptp2gps_conv_0:out_valid -> oran_tod_stack:i_ptp_master_tod_valid
	wire  [95:0] oran_ptp2gps_conv_0_gps_seconds_data;            // oran_ptp2gps_conv_0:gps_seconds -> oran_tod_stack:i_ptp_master_tod
	wire         master_tod_split_conduit_end_2_valid;            // master_tod_split:valid_conduit_out_2 -> oran_ptp2gps_conv_0:in_valid
	wire  [95:0] master_tod_split_conduit_end_2_data;             // master_tod_split:data_conduit_out_2 -> oran_ptp2gps_conv_0:ptp_seconds
	wire         tod_subsys_rst_100_out_reset_reset;              // tod_subsys_rst_100:out_reset_n -> [oran_tod_stack:i_reconfig_reset, port_8_tod_stack:i_reconfig_reset, rst_controller:reset_in0, tod_156_reset_controller_0:reset_in0]
	wire         tod_156_reset_controller_0_reset_out_reset;      // tod_156_reset_controller_0:reset_out -> oran_ptp2gps_conv_0:rst_tod_n
	wire         rst_controller_reset_out_reset;                  // rst_controller:reset_out -> [oran_tod_stack:i_ptp_master_tod_rst_n, port_8_tod_stack:i_ptp_master_tod_rst_n]

	master_tod_split master_tod_split (
		.data_conduit_in      (master_tod_split_conduit_end_data),     //   input,  width = 96,    conduit_end.data
		.valid_conduit_in     (master_tod_split_conduit_end_valid),    //   input,   width = 1,               .valid
		.data_conduit_out_1   (master_tod_split_conduit_end_1_data),   //  output,  width = 96,  conduit_end_1.data
		.valid_conduit_out_1  (master_tod_split_conduit_end_1_valid),  //  output,   width = 1,               .valid
		.data_conduit_out_2   (master_tod_split_conduit_end_2_data),   //  output,  width = 96,  conduit_end_2.data
		.valid_conduit_out_2  (master_tod_split_conduit_end_2_valid),  //  output,   width = 1,               .valid
		.data_conduit_out_3   (),                                      //  output,  width = 96,  conduit_end_3.data
		.valid_conduit_out_3  (),                                      //  output,   width = 1,               .valid
		.data_conduit_out_4   (),                                      //  output,  width = 96,  conduit_end_4.data
		.valid_conduit_out_4  (),                                      //  output,   width = 1,               .valid
		.data_conduit_out_5   (),                                      //  output,  width = 96,  conduit_end_5.data
		.valid_conduit_out_5  (),                                      //  output,   width = 1,               .valid
		.data_conduit_out_6   (),                                      //  output,  width = 96,  conduit_end_6.data
		.valid_conduit_out_6  (),                                      //  output,   width = 1,               .valid
		.data_conduit_out_7   (),                                      //  output,  width = 96,  conduit_end_7.data
		.valid_conduit_out_7  (),                                      //  output,   width = 1,               .valid
		.data_conduit_out_8   (),                                      //  output,  width = 96,  conduit_end_8.data
		.valid_conduit_out_8  (),                                      //  output,   width = 1,               .valid
		.data_conduit_out_9   (),                                      //  output,  width = 96,  conduit_end_9.data
		.valid_conduit_out_9  (),                                      //  output,   width = 1,               .valid
		.data_conduit_out_10  (master_tod_split_conduit_end_10_data),  //  output,  width = 96, conduit_end_10.data
		.valid_conduit_out_10 (master_tod_split_conduit_end_10_valid)  //  output,   width = 1,               .valid
	);

	oran_ptp2gps_conv_0 oran_ptp2gps_conv_0 (
		.rst_tod_n   (~tod_156_reset_controller_0_reset_out_reset), //   input,   width = 1,   rst_tod_n.reset_n
		.ptp_seconds (master_tod_split_conduit_end_2_data),         //   input,  width = 96, ptp_seconds.data
		.in_valid    (master_tod_split_conduit_end_2_valid),        //   input,   width = 1,            .valid
		.gps_seconds (oran_ptp2gps_conv_0_gps_seconds_data),        //  output,  width = 96, gps_seconds.data
		.out_valid   (oran_ptp2gps_conv_0_gps_seconds_valid),       //  output,   width = 1,            .valid
		.clk_tod     (tod_subsys_mtod_clk_out_clk_clk)              //   input,   width = 1,     clk_tod.clk
	);

	port_0_tod_stack_1 oran_tod_stack (
		.i_reconfig_clk              (tod_subsys_clk_100_out_clk_clk),                  //   input,   width = 1,          reconfig_clk.clk
		.i_reconfig_reset            (tod_subsys_rst_100_out_reset_reset),              //   input,   width = 1,       reconfig_resetn.reset_n
		.i_clk_tx_tod                (oran_tod_stack_tx_clk_clk),                       //   input,   width = 1,                tx_clk.clk
		.i_clk_rx_tod                (oran_tod_stack_rx_clk_clk),                       //   input,   width = 1,                rx_clk.clk
		.i_clk_master_tod            (tod_subsys_mtod_clk_out_clk_clk),                 //   input,   width = 1,              mtod_clk.clk
		.i_clk_todsync_sample        (oran_tod_stack_todsync_sample_clk_clk),           //   input,   width = 1,    todsync_sample_clk.clk
		.i_clk_todsync_sample_locked (todsync_sample_plllock_split_conduit_end_3_lock), //   input,   width = 1, todsync_sample_locked.lock
		.i_ptp_master_tod            (oran_ptp2gps_conv_0_gps_seconds_data),            //   input,  width = 96,  master_tod_interface.data
		.i_ptp_master_tod_valid      (oran_ptp2gps_conv_0_gps_seconds_valid),           //   input,   width = 1,                      .valid
		.ptp_tx_tod                  (oran_tod_stack_tx_tod_interface_tdata),           //  output,  width = 96,      tx_tod_interface.tdata
		.ptp_tx_tod_valid            (oran_tod_stack_tx_tod_interface_tvalid),          //  output,   width = 1,                      .tvalid
		.ptp_rx_tod                  (oran_tod_stack_rx_tod_interface_tdata),           //  output,  width = 96,      rx_tod_interface.tdata
		.ptp_rx_tod_valid            (oran_tod_stack_rx_tod_interface_tvalid),          //  output,   width = 1,                      .tvalid
		.i_tx_pll_locked             (oran_tod_stack_tx_pll_locked_lock),               //   input,   width = 1,         tx_pll_locked.lock
		.i_ptp_master_tod_rst_n      (~rst_controller_reset_out_reset)                  //   input,   width = 1,          mtod_reset_n.reset_n
	);

	port_0_tod_stack port_8_tod_stack (
		.i_reconfig_clk              (tod_subsys_clk_100_out_clk_clk),                  //   input,   width = 1,          reconfig_clk.clk
		.i_reconfig_reset            (tod_subsys_rst_100_out_reset_reset),              //   input,   width = 1,       reconfig_resetn.reset_n
		.i_clk_tx_tod                (port_8_tod_stack_tx_clk_clk),                     //   input,   width = 1,                tx_clk.clk
		.i_clk_rx_tod                (port_8_tod_stack_rx_clk_clk),                     //   input,   width = 1,                rx_clk.clk
		.i_clk_master_tod            (tod_subsys_mtod_clk_out_clk_clk),                 //   input,   width = 1,              mtod_clk.clk
		.i_clk_todsync_sample        (port_8_tod_stack_todsync_sample_clk_clk),         //   input,   width = 1,    todsync_sample_clk.clk
		.i_clk_todsync_sample_locked (todsync_sample_plllock_split_conduit_end_1_lock), //   input,   width = 1, todsync_sample_locked.lock
		.i_ptp_master_tod            (master_tod_split_conduit_end_1_data),             //   input,  width = 96,  master_tod_interface.data
		.i_ptp_master_tod_valid      (master_tod_split_conduit_end_1_valid),            //   input,   width = 1,                      .valid
		.ptp_tx_tod                  (port_8_tod_stack_tx_tod_interface_tdata),         //  output,  width = 96,      tx_tod_interface.tdata
		.ptp_tx_tod_valid            (port_8_tod_stack_tx_tod_interface_tvalid),        //  output,   width = 1,                      .tvalid
		.ptp_rx_tod                  (port_8_tod_stack_rx_tod_interface_tdata),         //  output,  width = 96,      rx_tod_interface.tdata
		.ptp_rx_tod_valid            (port_8_tod_stack_rx_tod_interface_tvalid),        //  output,   width = 1,                      .tvalid
		.i_tx_pll_locked             (port_8_tod_stack_tx_pll_locked_lock),             //   input,   width = 1,         tx_pll_locked.lock
		.i_ptp_master_tod_rst_n      (~rst_controller_reset_out_reset)                  //   input,   width = 1,          mtod_reset_n.reset_n
	);

	tod_156_reset_controller_0 tod_156_reset_controller_0 (
		.reset_in0 (~tod_subsys_rst_100_out_reset_reset),        //   input,  width = 1, reset_in0.reset
		.clk       (tod_subsys_mtod_clk_out_clk_clk),            //   input,  width = 1,       clk.clk
		.reset_out (tod_156_reset_controller_0_reset_out_reset)  //  output,  width = 1, reset_out.reset
	);

	tod_subsys_clk_100 tod_subsys_clk_100 (
		.in_clk  (tod_subsys_clk_100_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (tod_subsys_clk_100_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	tod_subsys_mtod_clk tod_subsys_mtod_clk (
		.in_clk  (tod_subsys_mtod_clk_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (tod_subsys_mtod_clk_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	tod_subsys_rst_100 tod_subsys_rst_100 (
		.clk         (tod_subsys_clk_100_out_clk_clk),      //   input,  width = 1,       clk.clk
		.in_reset_n  (tod_subsys_rst_100_in_reset_reset_n), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (tod_subsys_rst_100_out_reset_reset)   //  output,  width = 1, out_reset.reset_n
	);

	todsync_sample_plllock_split todsync_sample_plllock_split (
		.conduit_in     (todsync_sample_plllock_split_conduit_end_lock),   //   input,  width = 1,    conduit_end.lock
		.conduit_out_1  (todsync_sample_plllock_split_conduit_end_1_lock), //  output,  width = 1,  conduit_end_1.lock
		.conduit_out_2  (),                                                //  output,  width = 1,  conduit_end_2.lock
		.conduit_out_3  (todsync_sample_plllock_split_conduit_end_3_lock), //  output,  width = 1,  conduit_end_3.lock
		.conduit_out_4  (),                                                //  output,  width = 1,  conduit_end_4.lock
		.conduit_out_5  (),                                                //  output,  width = 1,  conduit_end_5.lock
		.conduit_out_6  (),                                                //  output,  width = 1,  conduit_end_6.lock
		.conduit_out_7  (),                                                //  output,  width = 1,  conduit_end_7.lock
		.conduit_out_8  (),                                                //  output,  width = 1,  conduit_end_8.lock
		.conduit_out_9  (),                                                //  output,  width = 1,  conduit_end_9.lock
		.conduit_out_10 (),                                                //  output,  width = 1, conduit_end_10.lock
		.conduit_out_11 (),                                                //  output,  width = 1, conduit_end_11.lock
		.conduit_out_12 (),                                                //  output,  width = 1, conduit_end_12.lock
		.conduit_out_13 (),                                                //  output,  width = 1, conduit_end_13.lock
		.conduit_out_14 (),                                                //  output,  width = 1, conduit_end_14.lock
		.conduit_out_15 (),                                                //  output,  width = 1, conduit_end_15.lock
		.conduit_out_16 (),                                                //  output,  width = 1, conduit_end_16.lock
		.conduit_out_17 (),                                                //  output,  width = 1, conduit_end_17.lock
		.conduit_out_18 (),                                                //  output,  width = 1, conduit_end_18.lock
		.conduit_out_19 (),                                                //  output,  width = 1, conduit_end_19.lock
		.conduit_out_20 ()                                                 //  output,  width = 1, conduit_end_20.lock
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~tod_subsys_rst_100_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (tod_subsys_mtod_clk_out_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      //  output,  width = 1, reset_out.reset
		.reset_req      (),                                    // (terminated),                       
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_in1      (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

endmodule
