/* ******************************************************************************************************************
 INTEL CONFIDENTIAL
 Copyright 2023 Intel Corporation All Rights Reserved.
 The source code contained or described herein and all documents related to the
 source code ("Material") are owned by Intel Corporation or its suppliers or
 licensors. Title to the Material remains with Intel Corporation or its
 suppliers and licensors. The Material may contain trade secrets and proprietary
 and confidential information of Intel Corporation and its suppliers and
 licensors, and is protected by worldwide copyright and trade secret laws and
 treaty provisions. No part of the Material may be used, copied, reproduced,
 modified, published, uploaded, posted, transmitted, distributed, or disclosed
 in any way without Intels prior express written permission.
 No license under any patent, copyright, trade secret or other intellectual
 property right is granted to or conferred upon you by disclosure or delivery
 of the Materials, either expressly, by implication, inducement, estoppel or
 otherwise. Any license under such intellectual property rights must be
 express and approved by Intel in writing.
 Unless otherwise agreed by Intel in writing, you may not remove or alter this
 notice or any other notice embedded in Materials by Intel or Intels suppliers
 or licensors in any way.
****************************************************************************************************************** */
`ifndef AVSTS_PKG_SV
`define AVSTS_PKG_SV

package  avsts_pkg;
  
  import uvm_pkg::*;
  `include "uvm_macros.svh"

   `include "../../avsts_uvc/items/avsts_item.sv"
   
   `include "../env/avsts_config.sv"
   `include "../env/avsts_sequencer.sv"
   `include "../env/avsts_monitor.sv"
   `include "../env/avsts_driver.sv"
   `include "../env/avsts_agent.sv"
   
   `include "../env/avsts_env.sv"
   
   `include "../sequences/avsts_sequences.sv"


endpackage :  avsts_pkg
`endif
