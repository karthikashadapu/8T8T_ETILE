// rst_ss.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module rst_ss (
		input  wire  dsp_rst_cntrl_reset_in0_reset,         //         dsp_rst_cntrl_reset_in0.reset
		input  wire  dsp_rst_cntrl_clk_clk,                 //               dsp_rst_cntrl_clk.clk
		output wire  dsp_rst_cntrl_reset_out_reset,         //         dsp_rst_cntrl_reset_out.reset
		input  wire  ecpri_rst_cntrl_reset_in0_reset,       //       ecpri_rst_cntrl_reset_in0.reset
		input  wire  ecpri_rst_cntrl_clk_clk,               //             ecpri_rst_cntrl_clk.clk
		output wire  ecpri_rst_cntrl_reset_out_reset,       //       ecpri_rst_cntrl_reset_out.reset
		input  wire  eth_rst_cntrl_reset_in0_reset,         //         eth_rst_cntrl_reset_in0.reset
		input  wire  eth_rst_cntrl_clk_clk,                 //               eth_rst_cntrl_clk.clk
		output wire  eth_rst_cntrl_reset_out_reset,         //         eth_rst_cntrl_reset_out.reset
		input  wire  reset_bridge_act_high_clk_clk,         //       reset_bridge_act_high_clk.clk
		input  wire  reset_bridge_act_high_in_reset_reset,  //  reset_bridge_act_high_in_reset.reset
		output wire  reset_bridge_act_high_out_reset_reset, // reset_bridge_act_high_out_reset.reset
		input  wire  rst_csr_clk_clk,                       //                     rst_csr_clk.clk
		input  wire  rst_csr_in_reset_reset_n,              //                rst_csr_in_reset.reset_n
		output wire  rst_csr_out_reset_reset_n,             //               rst_csr_out_reset.reset_n
		input  wire  reset_bridge_rec_rx_clk_clk,           //         reset_bridge_rec_rx_clk.clk
		input  wire  reset_bridge_rec_rx_in_reset_reset,    //    reset_bridge_rec_rx_in_reset.reset
		output wire  reset_bridge_rec_rx_out_reset_reset,   //   reset_bridge_rec_rx_out_reset.reset
		input  wire  reset_bridge_tx_div_clk_clk,           //         reset_bridge_tx_div_clk.clk
		input  wire  reset_bridge_tx_div_in_reset_reset,    //    reset_bridge_tx_div_in_reset.reset
		output wire  reset_bridge_tx_div_out_reset_reset    //   reset_bridge_tx_div_out_reset.reset
	);

	dsp_rst_cntrl dsp_rst_cntrl (
		.reset_in0 (dsp_rst_cntrl_reset_in0_reset), //   input,  width = 1, reset_in0.reset
		.clk       (dsp_rst_cntrl_clk_clk),         //   input,  width = 1,       clk.clk
		.reset_out (dsp_rst_cntrl_reset_out_reset)  //  output,  width = 1, reset_out.reset
	);

	ecpri_rst_cntrl ecpri_rst_cntrl (
		.reset_in0 (ecpri_rst_cntrl_reset_in0_reset), //   input,  width = 1, reset_in0.reset
		.clk       (ecpri_rst_cntrl_clk_clk),         //   input,  width = 1,       clk.clk
		.reset_out (ecpri_rst_cntrl_reset_out_reset)  //  output,  width = 1, reset_out.reset
	);

	eth_rst_cntrl eth_rst_cntrl (
		.reset_in0 (eth_rst_cntrl_reset_in0_reset), //   input,  width = 1, reset_in0.reset
		.clk       (eth_rst_cntrl_clk_clk),         //   input,  width = 1,       clk.clk
		.reset_out (eth_rst_cntrl_reset_out_reset)  //  output,  width = 1, reset_out.reset
	);

	reset_bridge_act_high reset_bridge_act_high (
		.clk       (reset_bridge_act_high_clk_clk),         //   input,  width = 1,       clk.clk
		.in_reset  (reset_bridge_act_high_in_reset_reset),  //   input,  width = 1,  in_reset.reset
		.out_reset (reset_bridge_act_high_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	rst_csr rst_csr (
		.clk         (rst_csr_clk_clk),           //   input,  width = 1,       clk.clk
		.in_reset_n  (rst_csr_in_reset_reset_n),  //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (rst_csr_out_reset_reset_n)  //  output,  width = 1, out_reset.reset_n
	);

	rst_ss_reset_bridge_rec_rx rst_ss_reset_bridge_rec_rx (
		.clk       (reset_bridge_rec_rx_clk_clk),         //   input,  width = 1,       clk.clk
		.in_reset  (reset_bridge_rec_rx_in_reset_reset),  //   input,  width = 1,  in_reset.reset
		.out_reset (reset_bridge_rec_rx_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	rst_ss_reset_bridge_tx_div rst_ss_reset_bridge_tx_div (
		.clk       (reset_bridge_tx_div_clk_clk),         //   input,  width = 1,       clk.clk
		.in_reset  (reset_bridge_tx_div_in_reset_reset),  //   input,  width = 1,  in_reset.reset
		.out_reset (reset_bridge_tx_div_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

endmodule
