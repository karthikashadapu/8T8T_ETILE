// lphy_ss_top.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module lphy_ss_top (
		input  wire         clk_csr_clk,                                    //                                    clk_csr.clk
		input  wire         clk_dsp_clk,                                    //                                    clk_dsp.clk
		input  wire         clk_xran_dl_clk,                                //                                clk_xran_dl.clk
		input  wire         clk_xran_ul_clk,                                //                                clk_xran_ul.clk
		output wire         pwr_mtr_h2f_bridge_s0_waitrequest,              //                      pwr_mtr_h2f_bridge_s0.waitrequest
		output wire [31:0]  pwr_mtr_h2f_bridge_s0_readdata,                 //                                           .readdata
		output wire         pwr_mtr_h2f_bridge_s0_readdatavalid,            //                                           .readdatavalid
		input  wire [0:0]   pwr_mtr_h2f_bridge_s0_burstcount,               //                                           .burstcount
		input  wire [31:0]  pwr_mtr_h2f_bridge_s0_writedata,                //                                           .writedata
		input  wire [16:0]  pwr_mtr_h2f_bridge_s0_address,                  //                                           .address
		input  wire         pwr_mtr_h2f_bridge_s0_write,                    //                                           .write
		input  wire         pwr_mtr_h2f_bridge_s0_read,                     //                                           .read
		input  wire [3:0]   pwr_mtr_h2f_bridge_s0_byteenable,               //                                           .byteenable
		input  wire         pwr_mtr_h2f_bridge_s0_debugaccess,              //                                           .debugaccess
		output wire         h2f_lw_bridge_s0_waitrequest,                   //                           h2f_lw_bridge_s0.waitrequest
		output wire [31:0]  h2f_lw_bridge_s0_readdata,                      //                                           .readdata
		output wire         h2f_lw_bridge_s0_readdatavalid,                 //                                           .readdatavalid
		input  wire [0:0]   h2f_lw_bridge_s0_burstcount,                    //                                           .burstcount
		input  wire [31:0]  h2f_lw_bridge_s0_writedata,                     //                                           .writedata
		input  wire [18:0]  h2f_lw_bridge_s0_address,                       //                                           .address
		input  wire         h2f_lw_bridge_s0_write,                         //                                           .write
		input  wire         h2f_lw_bridge_s0_read,                          //                                           .read
		input  wire [3:0]   h2f_lw_bridge_s0_byteenable,                    //                                           .byteenable
		input  wire         h2f_lw_bridge_s0_debugaccess,                   //                                           .debugaccess
		input  wire [16:0]  pb_mm_bridge_address,                           //                               pb_mm_bridge.address
		input  wire         pb_mm_bridge_chipselect,                        //                                           .chipselect
		input  wire         pb_mm_bridge_read,                              //                                           .read
		output wire [31:0]  pb_mm_bridge_readdata,                          //                                           .readdata
		input  wire         pb_mm_bridge_write,                             //                                           .write
		input  wire [31:0]  pb_mm_bridge_writedata,                         //                                           .writedata
		input  wire [3:0]   pb_mm_bridge_byteenable,                        //                                           .byteenable
		output wire         pb_mm_bridge_waitrequest,                       //                                           .waitrequest
		input  wire         xran_demapper_source_valid,                     //                       xran_demapper_source.valid
		input  wire [127:0] xran_demapper_source_data,                      //                                           .data
		input  wire         xran_demapper_source_endofpacket,               //                                           .endofpacket
		input  wire         xran_demapper_source_startofpacket,             //                                           .startofpacket
		output wire         xran_demapper_source_ready,                     //                                           .ready
		input  wire [15:0]  xran_demapper_source_channel,                   //                                           .channel
		output wire         ifft_source_l1_valid,                           //                             ifft_source_l1.valid
		output wire [31:0]  ifft_source_l1_data,                            //                                           .data
		output wire [7:0]   ifft_source_l1_channel,                         //                                           .channel
		output wire         ifft_source_l2_valid,                           //                             ifft_source_l2.valid
		output wire [31:0]  ifft_source_l2_data,                            //                                           .data
		output wire [7:0]   ifft_source_l2_channel,                         //                                           .channel
		output wire         coupling_pusch_avst_sink_l1_valid,              //                coupling_pusch_avst_sink_l1.valid
		output wire [31:0]  coupling_pusch_avst_sink_l1_data,               //                                           .data
		output wire [15:0]  coupling_pusch_avst_sink_l1_channel,            //                                           .channel
		output wire         coupling_pusch_avst_sink_l1_startofpacket,      //                                           .startofpacket
		output wire         coupling_pusch_avst_sink_l1_endofpacket,        //                                           .endofpacket
		output wire         coupling_pusch_avst_sink_l2_valid,              //                coupling_pusch_avst_sink_l2.valid
		output wire [31:0]  coupling_pusch_avst_sink_l2_data,               //                                           .data
		output wire [15:0]  coupling_pusch_avst_sink_l2_channel,            //                                           .channel
		output wire         coupling_pusch_avst_sink_l2_startofpacket,      //                                           .startofpacket
		output wire         coupling_pusch_avst_sink_l2_endofpacket,        //                                           .endofpacket
		output wire         coupling_prach_avst_sink_l1_valid,              //                coupling_prach_avst_sink_l1.valid
		output wire [31:0]  coupling_prach_avst_sink_l1_data,               //                                           .data
		output wire [15:0]  coupling_prach_avst_sink_l1_channel,            //                                           .channel
		output wire         coupling_prach_avst_sink_l1_startofpacket,      //                                           .startofpacket
		output wire         coupling_prach_avst_sink_l1_endofpacket,        //                                           .endofpacket
		output wire         coupling_prach_avst_sink_l2_valid,              //                coupling_prach_avst_sink_l2.valid
		output wire [31:0]  coupling_prach_avst_sink_l2_data,               //                                           .data
		output wire [15:0]  coupling_prach_avst_sink_l2_channel,            //                                           .channel
		output wire         coupling_prach_avst_sink_l2_startofpacket,      //                                           .startofpacket
		output wire         coupling_prach_avst_sink_l2_endofpacket,        //                                           .endofpacket
		input  wire         xran_demapper_cplane_source_valid,              //                xran_demapper_cplane_source.valid
		input  wire         xran_demapper_cplane_source_startofpacket,      //                                           .startofpacket
		input  wire         xran_demapper_cplane_source_endofpacket,        //                                           .endofpacket
		input  wire         pb_avst_sink_valid,                             //                               pb_avst_sink.valid
		input  wire [63:0]  pb_avst_sink_data,                              //                                           .data
		output wire         pb_avst_sink_ready,                             //                                           .ready
		output wire [7:0]   bw_confg_cc1_bw_config_cc1,                     //                               bw_confg_cc1.bw_config_cc1
		output wire [7:0]   bw_confg_cc2_bw_config_cc2,                     //                               bw_confg_cc2.bw_config_cc2
		output wire [55:0]  radio_config_status_radio_config_status,        //                        radio_config_status.radio_config_status
		output wire         short_long_prach_select_data,                   //                    short_long_prach_select.data
		input  wire [15:0]  rx_rtc_id_rx_rtc_id,                            //                                  rx_rtc_id.rx_rtc_id
		input  wire [15:0]  rx_u_axc_id_rx_u_axc_id,                        //                                rx_u_axc_id.rx_u_axc_id
		input  wire [15:0]  rx_rtc_id_dl_rx_rtc_id_dl,                      //                               rx_rtc_id_dl.rx_rtc_id_dl
		input  wire         lphy_ss_ul_sink_l1_valid,                       //                         lphy_ss_ul_sink_l1.valid
		input  wire [31:0]  lphy_ss_ul_sink_l1_data,                        //                                           .data
		input  wire [7:0]   lphy_ss_ul_sink_l1_channel,                     //                                           .channel
		input  wire         lphy_ss_ul_sink_l2_valid,                       //                         lphy_ss_ul_sink_l2.valid
		input  wire [31:0]  lphy_ss_ul_sink_l2_data,                        //                                           .data
		input  wire [7:0]   lphy_ss_ul_sink_l2_channel,                     //                                           .channel
		output wire         rst_soft_n_rst_soft_n,                          //                                 rst_soft_n.rst_soft_n
		output wire [31:0]  coupling_pusch_timing_ref_data,                 //                  coupling_pusch_timing_ref.data
		output wire [31:0]  coupling_prach_timing_ref_data,                 //                  coupling_prach_timing_ref.data
		input  wire [189:0] oran_rx_cplane_concat_data,                     //                      oran_rx_cplane_concat.data
		input  wire [67:0]  oran_rx_uplane_concat_data,                     //                      oran_rx_uplane_concat.data
		output wire         lphy_avst_selctd_cap_intf_valid,                //                  lphy_avst_selctd_cap_intf.valid
		output wire [31:0]  lphy_avst_selctd_cap_intf_data,                 //                                           .data
		output wire [2:0]   lphy_avst_selctd_cap_intf_channel,              //                                           .channel
		output wire         ul_start_pulse_latch_data,                      //                       ul_start_pulse_latch.data
		input  wire         frame_status_counter_reset_data,                //                 frame_status_counter_reset.data
		input  wire [31:0]  lphy_ss_top_interface_sel_data,                 //                  lphy_ss_top_interface_sel.data
		output wire         lphy_ss_top_dl_input_hfn_pulse_data,            //             lphy_ss_top_dl_input_hfn_pulse.data
		output wire         lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l1_irq, // lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l1.irq
		output wire         lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l2_irq, // lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l2.irq
		output wire         lphy_ss_top_pwr_mtr_fft_hist_done_intr_l1_irq,  //  lphy_ss_top_pwr_mtr_fft_hist_done_intr_l1.irq
		output wire         lphy_ss_top_pwr_mtr_fft_hist_done_intr_l2_irq,  //  lphy_ss_top_pwr_mtr_fft_hist_done_intr_l2.irq
		output wire         lphy_ss_top_duc_ddc_lpbk_en_data,               //                lphy_ss_top_duc_ddc_lpbk_en.data
		input  wire         reset_csr_reset,                                //                                  reset_csr.reset
		input  wire         reset_dsp_in_reset_n,                           //                               reset_dsp_in.reset_n
		input  wire         reset_xran_dl_reset_n,                          //                              reset_xran_dl.reset_n
		input  wire         reset_xran_ul_reset_n                           //                              reset_xran_ul.reset_n
	);

	wire         clk_xran_dl_out_clk_clk;                                                // clk_xran_dl:out_clk -> [lphy_ss_top:clk_eth_xran_dl, reset_xran_dl:clk]
	wire         clk_xran_ul_out_clk_clk;                                                // clk_xran_ul:out_clk -> [lphy_ss_top:clk_eth_xran_ul, reset_xran_ul:clk]
	wire         clk_csr_out_clk_clk;                                                    // clk_csr:out_clk -> [h2f_bridge:clk, h2f_lw_bridge:clk, lphy_ss_top:clk_csr, mm_interconnect_0:clk_csr_out_clk_clk, mm_interconnect_1:clk_csr_out_clk_clk, reset_csr:clk, rst_controller:clk]
	wire         clk_dsp_out_clk_clk;                                                    // clk_dsp:out_clk -> [lphy_ss_top:clk_dsp, reset_dsp:clk]
	wire         reset_csr_out_reset_reset;                                              // reset_csr:out_reset -> [h2f_bridge:reset, h2f_lw_bridge:reset, lphy_ss_top:rst_csr_n, rst_controller:reset_in0]
	wire         reset_dsp_out_reset_reset;                                              // reset_dsp:out_reset_n -> lphy_ss_top:rst_dsp_n
	wire         reset_xran_dl_out_reset_reset;                                          // reset_xran_dl:out_reset_n -> lphy_ss_top:rst_eth_xran_n_dl
	wire         reset_xran_ul_out_reset_reset;                                          // reset_xran_ul:out_reset_n -> lphy_ss_top:rst_eth_xran_n_ul
	wire         h2f_lw_bridge_m0_waitrequest;                                           // mm_interconnect_0:h2f_lw_bridge_m0_waitrequest -> h2f_lw_bridge:m0_waitrequest
	wire  [31:0] h2f_lw_bridge_m0_readdata;                                              // mm_interconnect_0:h2f_lw_bridge_m0_readdata -> h2f_lw_bridge:m0_readdata
	wire         h2f_lw_bridge_m0_debugaccess;                                           // h2f_lw_bridge:m0_debugaccess -> mm_interconnect_0:h2f_lw_bridge_m0_debugaccess
	wire  [18:0] h2f_lw_bridge_m0_address;                                               // h2f_lw_bridge:m0_address -> mm_interconnect_0:h2f_lw_bridge_m0_address
	wire         h2f_lw_bridge_m0_read;                                                  // h2f_lw_bridge:m0_read -> mm_interconnect_0:h2f_lw_bridge_m0_read
	wire   [3:0] h2f_lw_bridge_m0_byteenable;                                            // h2f_lw_bridge:m0_byteenable -> mm_interconnect_0:h2f_lw_bridge_m0_byteenable
	wire         h2f_lw_bridge_m0_readdatavalid;                                         // mm_interconnect_0:h2f_lw_bridge_m0_readdatavalid -> h2f_lw_bridge:m0_readdatavalid
	wire  [31:0] h2f_lw_bridge_m0_writedata;                                             // h2f_lw_bridge:m0_writedata -> mm_interconnect_0:h2f_lw_bridge_m0_writedata
	wire         h2f_lw_bridge_m0_write;                                                 // h2f_lw_bridge:m0_write -> mm_interconnect_0:h2f_lw_bridge_m0_write
	wire   [0:0] h2f_lw_bridge_m0_burstcount;                                            // h2f_lw_bridge:m0_burstcount -> mm_interconnect_0:h2f_lw_bridge_m0_burstcount
	wire  [31:0] mm_interconnect_0_lphy_ss_top_fft1_busin_readdata;                      // lphy_ss_top:fft1_busOut_readdata -> mm_interconnect_0:lphy_ss_top_fft1_busin_readdata
	wire         mm_interconnect_0_lphy_ss_top_fft1_busin_waitrequest;                   // lphy_ss_top:fft1_busOut_waitrequest -> mm_interconnect_0:lphy_ss_top_fft1_busin_waitrequest
	wire  [13:0] mm_interconnect_0_lphy_ss_top_fft1_busin_address;                       // mm_interconnect_0:lphy_ss_top_fft1_busin_address -> lphy_ss_top:fft1_busIn_address
	wire         mm_interconnect_0_lphy_ss_top_fft1_busin_read;                          // mm_interconnect_0:lphy_ss_top_fft1_busin_read -> lphy_ss_top:fft1_busIn_read
	wire         mm_interconnect_0_lphy_ss_top_fft1_busin_readdatavalid;                 // lphy_ss_top:fft1_busOut_readdatavalid -> mm_interconnect_0:lphy_ss_top_fft1_busin_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_fft1_busin_write;                         // mm_interconnect_0:lphy_ss_top_fft1_busin_write -> lphy_ss_top:fft1_busIn_write
	wire  [31:0] mm_interconnect_0_lphy_ss_top_fft1_busin_writedata;                     // mm_interconnect_0:lphy_ss_top_fft1_busin_writedata -> lphy_ss_top:fft1_busIn_writedata
	wire  [31:0] mm_interconnect_0_lphy_ss_top_fft2_busin_readdata;                      // lphy_ss_top:fft2_busOut_readdata -> mm_interconnect_0:lphy_ss_top_fft2_busin_readdata
	wire         mm_interconnect_0_lphy_ss_top_fft2_busin_waitrequest;                   // lphy_ss_top:fft2_busOut_waitrequest -> mm_interconnect_0:lphy_ss_top_fft2_busin_waitrequest
	wire  [13:0] mm_interconnect_0_lphy_ss_top_fft2_busin_address;                       // mm_interconnect_0:lphy_ss_top_fft2_busin_address -> lphy_ss_top:fft2_busIn_address
	wire         mm_interconnect_0_lphy_ss_top_fft2_busin_read;                          // mm_interconnect_0:lphy_ss_top_fft2_busin_read -> lphy_ss_top:fft2_busIn_read
	wire         mm_interconnect_0_lphy_ss_top_fft2_busin_readdatavalid;                 // lphy_ss_top:fft2_busOut_readdatavalid -> mm_interconnect_0:lphy_ss_top_fft2_busin_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_fft2_busin_write;                         // mm_interconnect_0:lphy_ss_top_fft2_busin_write -> lphy_ss_top:fft2_busIn_write
	wire  [31:0] mm_interconnect_0_lphy_ss_top_fft2_busin_writedata;                     // mm_interconnect_0:lphy_ss_top_fft2_busin_writedata -> lphy_ss_top:fft2_busIn_writedata
	wire  [31:0] mm_interconnect_0_lphy_ss_top_ifft1_busin_readdata;                     // lphy_ss_top:ifft1_busOut_readdata -> mm_interconnect_0:lphy_ss_top_ifft1_busin_readdata
	wire         mm_interconnect_0_lphy_ss_top_ifft1_busin_waitrequest;                  // lphy_ss_top:ifft1_busOut_waitrequest -> mm_interconnect_0:lphy_ss_top_ifft1_busin_waitrequest
	wire  [13:0] mm_interconnect_0_lphy_ss_top_ifft1_busin_address;                      // mm_interconnect_0:lphy_ss_top_ifft1_busin_address -> lphy_ss_top:ifft1_busIn_address
	wire         mm_interconnect_0_lphy_ss_top_ifft1_busin_read;                         // mm_interconnect_0:lphy_ss_top_ifft1_busin_read -> lphy_ss_top:ifft1_busIn_read
	wire         mm_interconnect_0_lphy_ss_top_ifft1_busin_readdatavalid;                // lphy_ss_top:ifft1_busOut_readdatavalid -> mm_interconnect_0:lphy_ss_top_ifft1_busin_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_ifft1_busin_write;                        // mm_interconnect_0:lphy_ss_top_ifft1_busin_write -> lphy_ss_top:ifft1_busIn_write
	wire  [31:0] mm_interconnect_0_lphy_ss_top_ifft1_busin_writedata;                    // mm_interconnect_0:lphy_ss_top_ifft1_busin_writedata -> lphy_ss_top:ifft1_busIn_writedata
	wire  [31:0] mm_interconnect_0_lphy_ss_top_ifft2_busin_readdata;                     // lphy_ss_top:ifft2_busOut_readdata -> mm_interconnect_0:lphy_ss_top_ifft2_busin_readdata
	wire         mm_interconnect_0_lphy_ss_top_ifft2_busin_waitrequest;                  // lphy_ss_top:ifft2_busOut_waitrequest -> mm_interconnect_0:lphy_ss_top_ifft2_busin_waitrequest
	wire  [13:0] mm_interconnect_0_lphy_ss_top_ifft2_busin_address;                      // mm_interconnect_0:lphy_ss_top_ifft2_busin_address -> lphy_ss_top:ifft2_busIn_address
	wire         mm_interconnect_0_lphy_ss_top_ifft2_busin_read;                         // mm_interconnect_0:lphy_ss_top_ifft2_busin_read -> lphy_ss_top:ifft2_busIn_read
	wire         mm_interconnect_0_lphy_ss_top_ifft2_busin_readdatavalid;                // lphy_ss_top:ifft2_busOut_readdatavalid -> mm_interconnect_0:lphy_ss_top_ifft2_busin_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_ifft2_busin_write;                        // mm_interconnect_0:lphy_ss_top_ifft2_busin_write -> lphy_ss_top:ifft2_busIn_write
	wire  [31:0] mm_interconnect_0_lphy_ss_top_ifft2_busin_writedata;                    // mm_interconnect_0:lphy_ss_top_ifft2_busin_writedata -> lphy_ss_top:ifft2_busIn_writedata
	wire  [31:0] mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_readdata;         // lphy_ss_top:long_prach_lw_bridge_readdata_l1 -> mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l1_readdata
	wire         mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_waitrequest;      // lphy_ss_top:long_prach_lw_bridge_waitrequest_l1 -> mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l1_waitrequest
	wire   [3:0] mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_address;          // mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l1_address -> lphy_ss_top:long_prach_lw_bridge_address_l1
	wire         mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_read;             // mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l1_read -> lphy_ss_top:long_prach_lw_bridge_read_l1
	wire         mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_readdatavalid;    // lphy_ss_top:long_prach_lw_bridge_readdatavalid_l1 -> mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l1_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_write;            // mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l1_write -> lphy_ss_top:long_prach_lw_bridge_write_l1
	wire  [31:0] mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_writedata;        // mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l1_writedata -> lphy_ss_top:long_prach_lw_bridge_writedata_l1
	wire  [31:0] mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_readdata;         // lphy_ss_top:long_prach_lw_bridge_readdata_l2 -> mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l2_readdata
	wire         mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_waitrequest;      // lphy_ss_top:long_prach_lw_bridge_waitrequest_l2 -> mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l2_waitrequest
	wire   [3:0] mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_address;          // mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l2_address -> lphy_ss_top:long_prach_lw_bridge_address_l2
	wire         mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_read;             // mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l2_read -> lphy_ss_top:long_prach_lw_bridge_read_l2
	wire         mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_readdatavalid;    // lphy_ss_top:long_prach_lw_bridge_readdatavalid_l2 -> mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l2_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_write;            // mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l2_write -> lphy_ss_top:long_prach_lw_bridge_write_l2
	wire  [31:0] mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_writedata;        // mm_interconnect_0:lphy_ss_top_long_prach_lw_bridge_l2_writedata -> lphy_ss_top:long_prach_lw_bridge_writedata_l2
	wire  [31:0] mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_readdata;              // lphy_ss_top:lphy_ss_config_csr_readdata -> mm_interconnect_0:lphy_ss_top_lphy_ss_config_csr_readdata
	wire         mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_waitrequest;           // lphy_ss_top:lphy_ss_config_csr_waitrequest -> mm_interconnect_0:lphy_ss_top_lphy_ss_config_csr_waitrequest
	wire   [7:0] mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_address;               // mm_interconnect_0:lphy_ss_top_lphy_ss_config_csr_address -> lphy_ss_top:lphy_ss_config_csr_address
	wire         mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_read;                  // mm_interconnect_0:lphy_ss_top_lphy_ss_config_csr_read -> lphy_ss_top:lphy_ss_config_csr_read
	wire         mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_readdatavalid;         // lphy_ss_top:lphy_ss_config_csr_readdatavalid -> mm_interconnect_0:lphy_ss_top_lphy_ss_config_csr_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_write;                 // mm_interconnect_0:lphy_ss_top_lphy_ss_config_csr_write -> lphy_ss_top:lphy_ss_config_csr_write
	wire  [31:0] mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_writedata;             // mm_interconnect_0:lphy_ss_top_lphy_ss_config_csr_writedata -> lphy_ss_top:lphy_ss_config_csr_writedata
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pb_ddr_csr_readdata;                      // lphy_ss_top:pb_ddr_csr_readdata -> mm_interconnect_0:lphy_ss_top_pb_ddr_csr_readdata
	wire   [3:0] mm_interconnect_0_lphy_ss_top_pb_ddr_csr_address;                       // mm_interconnect_0:lphy_ss_top_pb_ddr_csr_address -> lphy_ss_top:pb_ddr_csr_address
	wire         mm_interconnect_0_lphy_ss_top_pb_ddr_csr_write;                         // mm_interconnect_0:lphy_ss_top_pb_ddr_csr_write -> lphy_ss_top:pb_ddr_csr_write
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pb_ddr_csr_writedata;                     // mm_interconnect_0:lphy_ss_top_pb_ddr_csr_writedata -> lphy_ss_top:pb_ddr_csr_writedata
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdata;       // lphy_ss_top:pwr_mtr_fft_config_csr_readdata_l1 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdata
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_waitrequest;    // lphy_ss_top:pwr_mtr_fft_config_csr_waitrequest_l1 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l1_waitrequest
	wire   [3:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_address;        // mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l1_address -> lphy_ss_top:pwr_mtr_fft_config_csr_address_l1
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_read;           // mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l1_read -> lphy_ss_top:pwr_mtr_fft_config_csr_read_l1
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdatavalid;  // lphy_ss_top:pwr_mtr_fft_config_csr_readdatavalid_l1 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_write;          // mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l1_write -> lphy_ss_top:pwr_mtr_fft_config_csr_write_l1
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_writedata;      // mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l1_writedata -> lphy_ss_top:pwr_mtr_fft_config_csr_writedata_l1
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdata;       // lphy_ss_top:pwr_mtr_fft_config_csr_readdata_l2 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdata
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_waitrequest;    // lphy_ss_top:pwr_mtr_fft_config_csr_waitrequest_l2 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l2_waitrequest
	wire   [3:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_address;        // mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l2_address -> lphy_ss_top:pwr_mtr_fft_config_csr_address_l2
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_read;           // mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l2_read -> lphy_ss_top:pwr_mtr_fft_config_csr_read_l2
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdatavalid;  // lphy_ss_top:pwr_mtr_fft_config_csr_readdatavalid_l2 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_write;          // mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l2_write -> lphy_ss_top:pwr_mtr_fft_config_csr_write_l2
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_writedata;      // mm_interconnect_0:lphy_ss_top_pwr_mtr_fft_config_csr_l2_writedata -> lphy_ss_top:pwr_mtr_fft_config_csr_writedata_l2
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdata;      // lphy_ss_top:pwr_mtr_ifft_config_csr_readdata_l1 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdata
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_waitrequest;   // lphy_ss_top:pwr_mtr_ifft_config_csr_waitrequest_l1 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l1_waitrequest
	wire   [3:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_address;       // mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l1_address -> lphy_ss_top:pwr_mtr_ifft_config_csr_address_l1
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_read;          // mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l1_read -> lphy_ss_top:pwr_mtr_ifft_config_csr_read_l1
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdatavalid; // lphy_ss_top:pwr_mtr_ifft_config_csr_readdatavalid_l1 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_write;         // mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l1_write -> lphy_ss_top:pwr_mtr_ifft_config_csr_write_l1
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_writedata;     // mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l1_writedata -> lphy_ss_top:pwr_mtr_ifft_config_csr_writedata_l1
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdata;      // lphy_ss_top:pwr_mtr_ifft_config_csr_readdata_l2 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdata
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_waitrequest;   // lphy_ss_top:pwr_mtr_ifft_config_csr_waitrequest_l2 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l2_waitrequest
	wire   [3:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_address;       // mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l2_address -> lphy_ss_top:pwr_mtr_ifft_config_csr_address_l2
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_read;          // mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l2_read -> lphy_ss_top:pwr_mtr_ifft_config_csr_read_l2
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdatavalid; // lphy_ss_top:pwr_mtr_ifft_config_csr_readdatavalid_l2 -> mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_write;         // mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l2_write -> lphy_ss_top:pwr_mtr_ifft_config_csr_write_l2
	wire  [31:0] mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_writedata;     // mm_interconnect_0:lphy_ss_top_pwr_mtr_ifft_config_csr_l2_writedata -> lphy_ss_top:pwr_mtr_ifft_config_csr_writedata_l2
	wire  [31:0] mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_readdata;        // lphy_ss_top:short_prach1_busOut_readdata -> mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l1_readdata
	wire         mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_waitrequest;     // lphy_ss_top:short_prach1_busOut_waitrequest -> mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l1_waitrequest
	wire   [9:0] mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_address;         // mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l1_address -> lphy_ss_top:short_prach1_busIn_address
	wire         mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_read;            // mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l1_read -> lphy_ss_top:short_prach1_busIn_read
	wire         mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_readdatavalid;   // lphy_ss_top:short_prach1_busOut_readdatavalid -> mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l1_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_write;           // mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l1_write -> lphy_ss_top:short_prach1_busIn_write
	wire  [31:0] mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_writedata;       // mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l1_writedata -> lphy_ss_top:short_prach1_busIn_writedata
	wire  [31:0] mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_readdata;        // lphy_ss_top:short_prach2_busOut_readdata -> mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l2_readdata
	wire         mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_waitrequest;     // lphy_ss_top:short_prach2_busOut_waitrequest -> mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l2_waitrequest
	wire   [9:0] mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_address;         // mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l2_address -> lphy_ss_top:short_prach2_busIn_address
	wire         mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_read;            // mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l2_read -> lphy_ss_top:short_prach2_busIn_read
	wire         mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_readdatavalid;   // lphy_ss_top:short_prach2_busOut_readdatavalid -> mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l2_readdatavalid
	wire         mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_write;           // mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l2_write -> lphy_ss_top:short_prach2_busIn_write
	wire  [31:0] mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_writedata;       // mm_interconnect_0:lphy_ss_top_short_prach_lw_bridge_l2_writedata -> lphy_ss_top:short_prach2_busIn_writedata
	wire         h2f_bridge_m0_waitrequest;                                              // mm_interconnect_1:h2f_bridge_m0_waitrequest -> h2f_bridge:m0_waitrequest
	wire  [31:0] h2f_bridge_m0_readdata;                                                 // mm_interconnect_1:h2f_bridge_m0_readdata -> h2f_bridge:m0_readdata
	wire         h2f_bridge_m0_debugaccess;                                              // h2f_bridge:m0_debugaccess -> mm_interconnect_1:h2f_bridge_m0_debugaccess
	wire  [16:0] h2f_bridge_m0_address;                                                  // h2f_bridge:m0_address -> mm_interconnect_1:h2f_bridge_m0_address
	wire         h2f_bridge_m0_read;                                                     // h2f_bridge:m0_read -> mm_interconnect_1:h2f_bridge_m0_read
	wire   [3:0] h2f_bridge_m0_byteenable;                                               // h2f_bridge:m0_byteenable -> mm_interconnect_1:h2f_bridge_m0_byteenable
	wire         h2f_bridge_m0_readdatavalid;                                            // mm_interconnect_1:h2f_bridge_m0_readdatavalid -> h2f_bridge:m0_readdatavalid
	wire  [31:0] h2f_bridge_m0_writedata;                                                // h2f_bridge:m0_writedata -> mm_interconnect_1:h2f_bridge_m0_writedata
	wire         h2f_bridge_m0_write;                                                    // h2f_bridge:m0_write -> mm_interconnect_1:h2f_bridge_m0_write
	wire   [0:0] h2f_bridge_m0_burstcount;                                               // h2f_bridge:m0_burstcount -> mm_interconnect_1:h2f_bridge_m0_burstcount
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_chipselect;      // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_chipselect -> lphy_ss_top:pm_fft_hist_mm_bridge_chipselect_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdata;        // lphy_ss_top:pm_fft_hist_mm_bridge_readdata_l1 -> mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_waitrequest;     // lphy_ss_top:pm_fft_hist_mm_bridge_waitrequest_l1 -> mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_waitrequest
	wire  [11:0] mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_address;         // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_address -> lphy_ss_top:pm_fft_hist_mm_bridge_address_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_read;            // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_read -> lphy_ss_top:pm_fft_hist_mm_bridge_read_l1
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_byteenable;      // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_byteenable -> lphy_ss_top:pm_fft_hist_mm_bridge_byteenable_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdatavalid;   // lphy_ss_top:pm_fft_hist_mm_bridge_readdatavalid_l1 -> mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdatavalid
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_write;           // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_write -> lphy_ss_top:pm_fft_hist_mm_bridge_write_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_writedata;       // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l1_writedata -> lphy_ss_top:pm_fft_hist_mm_bridge_writedata_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_chipselect;      // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_chipselect -> lphy_ss_top:pm_fft_hist_mm_bridge_chipselect_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdata;        // lphy_ss_top:pm_fft_hist_mm_bridge_readdata_l2 -> mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_waitrequest;     // lphy_ss_top:pm_fft_hist_mm_bridge_waitrequest_l2 -> mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_waitrequest
	wire  [11:0] mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_address;         // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_address -> lphy_ss_top:pm_fft_hist_mm_bridge_address_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_read;            // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_read -> lphy_ss_top:pm_fft_hist_mm_bridge_read_l2
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_byteenable;      // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_byteenable -> lphy_ss_top:pm_fft_hist_mm_bridge_byteenable_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdatavalid;   // lphy_ss_top:pm_fft_hist_mm_bridge_readdatavalid_l2 -> mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdatavalid
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_write;           // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_write -> lphy_ss_top:pm_fft_hist_mm_bridge_write_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_writedata;       // mm_interconnect_1:lphy_ss_top_pm_fft_hist_mm_bridge_l2_writedata -> lphy_ss_top:pm_fft_hist_mm_bridge_writedata_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_chipselect;   // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l1_chipselect -> lphy_ss_top:pm_fft_threash_mm_bridge_chipselect_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_readdata;     // lphy_ss_top:pm_fft_threash_mm_bridge_readdata_l1 -> mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l1_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_waitrequest;  // lphy_ss_top:pm_fft_threash_mm_bridge_waitrequest_l1 -> mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l1_waitrequest
	wire   [5:0] mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_address;      // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l1_address -> lphy_ss_top:pm_fft_threash_mm_bridge_address_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_read;         // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l1_read -> lphy_ss_top:pm_fft_threash_mm_bridge_read_l1
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_byteenable;   // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l1_byteenable -> lphy_ss_top:pm_fft_threash_mm_bridge_byteenable_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_write;        // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l1_write -> lphy_ss_top:pm_fft_threash_mm_bridge_write_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_writedata;    // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l1_writedata -> lphy_ss_top:pm_fft_threash_mm_bridge_writedata_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_chipselect;   // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l2_chipselect -> lphy_ss_top:pm_fft_threash_mm_bridge_chipselect_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_readdata;     // lphy_ss_top:pm_fft_threash_mm_bridge_readdata_l2 -> mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l2_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_waitrequest;  // lphy_ss_top:pm_fft_threash_mm_bridge_waitrequest_l2 -> mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l2_waitrequest
	wire   [5:0] mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_address;      // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l2_address -> lphy_ss_top:pm_fft_threash_mm_bridge_address_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_read;         // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l2_read -> lphy_ss_top:pm_fft_threash_mm_bridge_read_l2
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_byteenable;   // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l2_byteenable -> lphy_ss_top:pm_fft_threash_mm_bridge_byteenable_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_write;        // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l2_write -> lphy_ss_top:pm_fft_threash_mm_bridge_write_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_writedata;    // mm_interconnect_1:lphy_ss_top_pm_fft_threash_mm_bridge_l2_writedata -> lphy_ss_top:pm_fft_threash_mm_bridge_writedata_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_chipselect;     // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_chipselect -> lphy_ss_top:pm_ifft_hist_mm_bridge_chipselect_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdata;       // lphy_ss_top:pm_ifft_hist_mm_bridge_readdata_l1 -> mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_waitrequest;    // lphy_ss_top:pm_ifft_hist_mm_bridge_waitrequest_l1 -> mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_waitrequest
	wire  [11:0] mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_address;        // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_address -> lphy_ss_top:pm_ifft_hist_mm_bridge_address_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_read;           // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_read -> lphy_ss_top:pm_ifft_hist_mm_bridge_read_l1
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_byteenable;     // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_byteenable -> lphy_ss_top:pm_ifft_hist_mm_bridge_byteenable_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdatavalid;  // lphy_ss_top:pm_ifft_hist_mm_bridge_readdatavalid_l1 -> mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdatavalid
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_write;          // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_write -> lphy_ss_top:pm_ifft_hist_mm_bridge_write_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_writedata;      // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l1_writedata -> lphy_ss_top:pm_ifft_hist_mm_bridge_writedata_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_chipselect;     // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_chipselect -> lphy_ss_top:pm_ifft_hist_mm_bridge_chipselect_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdata;       // lphy_ss_top:pm_ifft_hist_mm_bridge_readdata_l2 -> mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_waitrequest;    // lphy_ss_top:pm_ifft_hist_mm_bridge_waitrequest_l2 -> mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_waitrequest
	wire  [11:0] mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_address;        // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_address -> lphy_ss_top:pm_ifft_hist_mm_bridge_address_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_read;           // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_read -> lphy_ss_top:pm_ifft_hist_mm_bridge_read_l2
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_byteenable;     // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_byteenable -> lphy_ss_top:pm_ifft_hist_mm_bridge_byteenable_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdatavalid;  // lphy_ss_top:pm_ifft_hist_mm_bridge_readdatavalid_l2 -> mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdatavalid
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_write;          // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_write -> lphy_ss_top:pm_ifft_hist_mm_bridge_write_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_writedata;      // mm_interconnect_1:lphy_ss_top_pm_ifft_hist_mm_bridge_l2_writedata -> lphy_ss_top:pm_ifft_hist_mm_bridge_writedata_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_chipselect;  // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l1_chipselect -> lphy_ss_top:pm_ifft_threash_mm_bridge_chipselect_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_readdata;    // lphy_ss_top:pm_ifft_threash_mm_bridge_readdata_l1 -> mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l1_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_waitrequest; // lphy_ss_top:pm_ifft_threash_mm_bridge_waitrequest_l1 -> mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l1_waitrequest
	wire   [5:0] mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_address;     // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l1_address -> lphy_ss_top:pm_ifft_threash_mm_bridge_address_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_read;        // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l1_read -> lphy_ss_top:pm_ifft_threash_mm_bridge_read_l1
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_byteenable;  // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l1_byteenable -> lphy_ss_top:pm_ifft_threash_mm_bridge_byteenable_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_write;       // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l1_write -> lphy_ss_top:pm_ifft_threash_mm_bridge_write_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_writedata;   // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l1_writedata -> lphy_ss_top:pm_ifft_threash_mm_bridge_writedata_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_chipselect;  // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l2_chipselect -> lphy_ss_top:pm_ifft_threash_mm_bridge_chipselect_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_readdata;    // lphy_ss_top:pm_ifft_threash_mm_bridge_readdata_l2 -> mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l2_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_waitrequest; // lphy_ss_top:pm_ifft_threash_mm_bridge_waitrequest_l2 -> mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l2_waitrequest
	wire   [5:0] mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_address;     // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l2_address -> lphy_ss_top:pm_ifft_threash_mm_bridge_address_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_read;        // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l2_read -> lphy_ss_top:pm_ifft_threash_mm_bridge_read_l2
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_byteenable;  // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l2_byteenable -> lphy_ss_top:pm_ifft_threash_mm_bridge_byteenable_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_write;       // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l2_write -> lphy_ss_top:pm_ifft_threash_mm_bridge_write_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_writedata;   // mm_interconnect_1:lphy_ss_top_pm_ifft_threash_mm_bridge_l2_writedata -> lphy_ss_top:pm_ifft_threash_mm_bridge_writedata_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_chipselect;      // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_chipselect -> lphy_ss_top:pm_stat_fft_mm_bridge_chipselect_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdata;        // lphy_ss_top:pm_stat_fft_mm_bridge_readdata_l1 -> mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_waitrequest;     // lphy_ss_top:pm_stat_fft_mm_bridge_waitrequest_l1 -> mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_waitrequest
	wire   [9:0] mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_address;         // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_address -> lphy_ss_top:pm_stat_fft_mm_bridge_address_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_read;            // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_read -> lphy_ss_top:pm_stat_fft_mm_bridge_read_l1
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_byteenable;      // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_byteenable -> lphy_ss_top:pm_stat_fft_mm_bridge_byteenable_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdatavalid;   // lphy_ss_top:pm_stat_fft_mm_bridge_readdatavalid_l1 -> mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdatavalid
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_write;           // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_write -> lphy_ss_top:pm_stat_fft_mm_bridge_write_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_writedata;       // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l1_writedata -> lphy_ss_top:pm_stat_fft_mm_bridge_writedata_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_chipselect;      // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_chipselect -> lphy_ss_top:pm_stat_fft_mm_bridge_chipselect_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdata;        // lphy_ss_top:pm_stat_fft_mm_bridge_readdata_l2 -> mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_waitrequest;     // lphy_ss_top:pm_stat_fft_mm_bridge_waitrequest_l2 -> mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_waitrequest
	wire   [9:0] mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_address;         // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_address -> lphy_ss_top:pm_stat_fft_mm_bridge_address_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_read;            // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_read -> lphy_ss_top:pm_stat_fft_mm_bridge_read_l2
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_byteenable;      // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_byteenable -> lphy_ss_top:pm_stat_fft_mm_bridge_byteenable_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdatavalid;   // lphy_ss_top:pm_stat_fft_mm_bridge_readdatavalid_l2 -> mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdatavalid
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_write;           // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_write -> lphy_ss_top:pm_stat_fft_mm_bridge_write_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_writedata;       // mm_interconnect_1:lphy_ss_top_pm_stat_fft_mm_bridge_l2_writedata -> lphy_ss_top:pm_stat_fft_mm_bridge_writedata_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_chipselect;     // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_chipselect -> lphy_ss_top:pm_stat_ifft_mm_bridge_chipselect_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdata;       // lphy_ss_top:pm_stat_ifft_mm_bridge_readdata_l1 -> mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_waitrequest;    // lphy_ss_top:pm_stat_ifft_mm_bridge_waitrequest_l1 -> mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_waitrequest
	wire   [9:0] mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_address;        // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_address -> lphy_ss_top:pm_stat_ifft_mm_bridge_address_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_read;           // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_read -> lphy_ss_top:pm_stat_ifft_mm_bridge_read_l1
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_byteenable;     // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_byteenable -> lphy_ss_top:pm_stat_ifft_mm_bridge_byteenable_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdatavalid;  // lphy_ss_top:pm_stat_ifft_mm_bridge_readdatavalid_l1 -> mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdatavalid
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_write;          // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_write -> lphy_ss_top:pm_stat_ifft_mm_bridge_write_l1
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_writedata;      // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l1_writedata -> lphy_ss_top:pm_stat_ifft_mm_bridge_writedata_l1
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_chipselect;     // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_chipselect -> lphy_ss_top:pm_stat_ifft_mm_bridge_chipselect_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdata;       // lphy_ss_top:pm_stat_ifft_mm_bridge_readdata_l2 -> mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdata
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_waitrequest;    // lphy_ss_top:pm_stat_ifft_mm_bridge_waitrequest_l2 -> mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_waitrequest
	wire   [9:0] mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_address;        // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_address -> lphy_ss_top:pm_stat_ifft_mm_bridge_address_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_read;           // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_read -> lphy_ss_top:pm_stat_ifft_mm_bridge_read_l2
	wire   [3:0] mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_byteenable;     // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_byteenable -> lphy_ss_top:pm_stat_ifft_mm_bridge_byteenable_l2
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdatavalid;  // lphy_ss_top:pm_stat_ifft_mm_bridge_readdatavalid_l2 -> mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdatavalid
	wire         mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_write;          // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_write -> lphy_ss_top:pm_stat_ifft_mm_bridge_write_l2
	wire  [31:0] mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_writedata;      // mm_interconnect_1:lphy_ss_top_pm_stat_ifft_mm_bridge_l2_writedata -> lphy_ss_top:pm_stat_ifft_mm_bridge_writedata_l2
	wire         rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [mm_interconnect_0:h2f_lw_bridge_m0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:h2f_lw_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:h2f_bridge_m0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:h2f_bridge_reset_reset_bridge_in_reset_reset]

	lphy_ss_clk_csr clk_csr (
		.in_clk  (clk_csr_clk),         //   input,  width = 1,  in_clk.clk
		.out_clk (clk_csr_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	lphy_ss_clk_dsp clk_dsp (
		.in_clk  (clk_dsp_clk),         //   input,  width = 1,  in_clk.clk
		.out_clk (clk_dsp_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	lphy_ss_clk_xran_dl clk_xran_dl (
		.in_clk  (clk_xran_dl_clk),         //   input,  width = 1,  in_clk.clk
		.out_clk (clk_xran_dl_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	lphy_ss_clk_xran_ul clk_xran_ul (
		.in_clk  (clk_xran_ul_clk),         //   input,  width = 1,  in_clk.clk
		.out_clk (clk_xran_ul_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	lphy_ss_top_h2f_bridge h2f_bridge (
		.clk              (clk_csr_out_clk_clk),                 //   input,   width = 1,   clk.clk
		.reset            (reset_csr_out_reset_reset),           //   input,   width = 1, reset.reset
		.s0_waitrequest   (pwr_mtr_h2f_bridge_s0_waitrequest),   //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (pwr_mtr_h2f_bridge_s0_readdata),      //  output,  width = 32,      .readdata
		.s0_readdatavalid (pwr_mtr_h2f_bridge_s0_readdatavalid), //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (pwr_mtr_h2f_bridge_s0_burstcount),    //   input,   width = 1,      .burstcount
		.s0_writedata     (pwr_mtr_h2f_bridge_s0_writedata),     //   input,  width = 32,      .writedata
		.s0_address       (pwr_mtr_h2f_bridge_s0_address),       //   input,  width = 17,      .address
		.s0_write         (pwr_mtr_h2f_bridge_s0_write),         //   input,   width = 1,      .write
		.s0_read          (pwr_mtr_h2f_bridge_s0_read),          //   input,   width = 1,      .read
		.s0_byteenable    (pwr_mtr_h2f_bridge_s0_byteenable),    //   input,   width = 4,      .byteenable
		.s0_debugaccess   (pwr_mtr_h2f_bridge_s0_debugaccess),   //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (h2f_bridge_m0_waitrequest),           //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (h2f_bridge_m0_readdata),              //   input,  width = 32,      .readdata
		.m0_readdatavalid (h2f_bridge_m0_readdatavalid),         //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (h2f_bridge_m0_burstcount),            //  output,   width = 1,      .burstcount
		.m0_writedata     (h2f_bridge_m0_writedata),             //  output,  width = 32,      .writedata
		.m0_address       (h2f_bridge_m0_address),               //  output,  width = 17,      .address
		.m0_write         (h2f_bridge_m0_write),                 //  output,   width = 1,      .write
		.m0_read          (h2f_bridge_m0_read),                  //  output,   width = 1,      .read
		.m0_byteenable    (h2f_bridge_m0_byteenable),            //  output,   width = 4,      .byteenable
		.m0_debugaccess   (h2f_bridge_m0_debugaccess)            //  output,   width = 1,      .debugaccess
	);

	lphy_ss_top_mm_bridge_0 h2f_lw_bridge (
		.clk              (clk_csr_out_clk_clk),            //   input,   width = 1,   clk.clk
		.reset            (reset_csr_out_reset_reset),      //   input,   width = 1, reset.reset
		.s0_waitrequest   (h2f_lw_bridge_s0_waitrequest),   //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (h2f_lw_bridge_s0_readdata),      //  output,  width = 32,      .readdata
		.s0_readdatavalid (h2f_lw_bridge_s0_readdatavalid), //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (h2f_lw_bridge_s0_burstcount),    //   input,   width = 1,      .burstcount
		.s0_writedata     (h2f_lw_bridge_s0_writedata),     //   input,  width = 32,      .writedata
		.s0_address       (h2f_lw_bridge_s0_address),       //   input,  width = 19,      .address
		.s0_write         (h2f_lw_bridge_s0_write),         //   input,   width = 1,      .write
		.s0_read          (h2f_lw_bridge_s0_read),          //   input,   width = 1,      .read
		.s0_byteenable    (h2f_lw_bridge_s0_byteenable),    //   input,   width = 4,      .byteenable
		.s0_debugaccess   (h2f_lw_bridge_s0_debugaccess),   //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (h2f_lw_bridge_m0_waitrequest),   //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (h2f_lw_bridge_m0_readdata),      //   input,  width = 32,      .readdata
		.m0_readdatavalid (h2f_lw_bridge_m0_readdatavalid), //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (h2f_lw_bridge_m0_burstcount),    //  output,   width = 1,      .burstcount
		.m0_writedata     (h2f_lw_bridge_m0_writedata),     //  output,  width = 32,      .writedata
		.m0_address       (h2f_lw_bridge_m0_address),       //  output,  width = 19,      .address
		.m0_write         (h2f_lw_bridge_m0_write),         //  output,   width = 1,      .write
		.m0_read          (h2f_lw_bridge_m0_read),          //  output,   width = 1,      .read
		.m0_byteenable    (h2f_lw_bridge_m0_byteenable),    //  output,   width = 4,      .byteenable
		.m0_debugaccess   (h2f_lw_bridge_m0_debugaccess)    //  output,   width = 1,      .debugaccess
	);

	lphy_ss_lphy_ss_top lphy_ss_top (
		.ifft1_busIn_writedata                    (mm_interconnect_0_lphy_ss_top_ifft1_busin_writedata),                    //   input,   width = 32,                    ifft1_busin.writedata
		.ifft1_busIn_address                      (mm_interconnect_0_lphy_ss_top_ifft1_busin_address),                      //   input,   width = 14,                               .address
		.ifft1_busIn_write                        (mm_interconnect_0_lphy_ss_top_ifft1_busin_write),                        //   input,    width = 1,                               .write
		.ifft1_busIn_read                         (mm_interconnect_0_lphy_ss_top_ifft1_busin_read),                         //   input,    width = 1,                               .read
		.ifft1_busOut_readdatavalid               (mm_interconnect_0_lphy_ss_top_ifft1_busin_readdatavalid),                //  output,    width = 1,                               .readdatavalid
		.ifft1_busOut_readdata                    (mm_interconnect_0_lphy_ss_top_ifft1_busin_readdata),                     //  output,   width = 32,                               .readdata
		.ifft1_busOut_waitrequest                 (mm_interconnect_0_lphy_ss_top_ifft1_busin_waitrequest),                  //  output,    width = 1,                               .waitrequest
		.ifft2_busIn_writedata                    (mm_interconnect_0_lphy_ss_top_ifft2_busin_writedata),                    //   input,   width = 32,                    ifft2_busin.writedata
		.ifft2_busIn_address                      (mm_interconnect_0_lphy_ss_top_ifft2_busin_address),                      //   input,   width = 14,                               .address
		.ifft2_busIn_write                        (mm_interconnect_0_lphy_ss_top_ifft2_busin_write),                        //   input,    width = 1,                               .write
		.ifft2_busIn_read                         (mm_interconnect_0_lphy_ss_top_ifft2_busin_read),                         //   input,    width = 1,                               .read
		.ifft2_busOut_readdatavalid               (mm_interconnect_0_lphy_ss_top_ifft2_busin_readdatavalid),                //  output,    width = 1,                               .readdatavalid
		.ifft2_busOut_readdata                    (mm_interconnect_0_lphy_ss_top_ifft2_busin_readdata),                     //  output,   width = 32,                               .readdata
		.ifft2_busOut_waitrequest                 (mm_interconnect_0_lphy_ss_top_ifft2_busin_waitrequest),                  //  output,    width = 1,                               .waitrequest
		.fft1_busIn_writedata                     (mm_interconnect_0_lphy_ss_top_fft1_busin_writedata),                     //   input,   width = 32,                     fft1_busin.writedata
		.fft1_busIn_address                       (mm_interconnect_0_lphy_ss_top_fft1_busin_address),                       //   input,   width = 14,                               .address
		.fft1_busIn_write                         (mm_interconnect_0_lphy_ss_top_fft1_busin_write),                         //   input,    width = 1,                               .write
		.fft1_busIn_read                          (mm_interconnect_0_lphy_ss_top_fft1_busin_read),                          //   input,    width = 1,                               .read
		.fft1_busOut_readdatavalid                (mm_interconnect_0_lphy_ss_top_fft1_busin_readdatavalid),                 //  output,    width = 1,                               .readdatavalid
		.fft1_busOut_readdata                     (mm_interconnect_0_lphy_ss_top_fft1_busin_readdata),                      //  output,   width = 32,                               .readdata
		.fft1_busOut_waitrequest                  (mm_interconnect_0_lphy_ss_top_fft1_busin_waitrequest),                   //  output,    width = 1,                               .waitrequest
		.fft2_busIn_writedata                     (mm_interconnect_0_lphy_ss_top_fft2_busin_writedata),                     //   input,   width = 32,                     fft2_busin.writedata
		.fft2_busIn_address                       (mm_interconnect_0_lphy_ss_top_fft2_busin_address),                       //   input,   width = 14,                               .address
		.fft2_busIn_write                         (mm_interconnect_0_lphy_ss_top_fft2_busin_write),                         //   input,    width = 1,                               .write
		.fft2_busIn_read                          (mm_interconnect_0_lphy_ss_top_fft2_busin_read),                          //   input,    width = 1,                               .read
		.fft2_busOut_readdatavalid                (mm_interconnect_0_lphy_ss_top_fft2_busin_readdatavalid),                 //  output,    width = 1,                               .readdatavalid
		.fft2_busOut_readdata                     (mm_interconnect_0_lphy_ss_top_fft2_busin_readdata),                      //  output,   width = 32,                               .readdata
		.fft2_busOut_waitrequest                  (mm_interconnect_0_lphy_ss_top_fft2_busin_waitrequest),                   //  output,    width = 1,                               .waitrequest
		.pb_ddr_csr_address                       (mm_interconnect_0_lphy_ss_top_pb_ddr_csr_address),                       //   input,    width = 4,                     pb_ddr_csr.address
		.pb_ddr_csr_write                         (mm_interconnect_0_lphy_ss_top_pb_ddr_csr_write),                         //   input,    width = 1,                               .write
		.pb_ddr_csr_writedata                     (mm_interconnect_0_lphy_ss_top_pb_ddr_csr_writedata),                     //   input,   width = 32,                               .writedata
		.pb_ddr_csr_readdata                      (mm_interconnect_0_lphy_ss_top_pb_ddr_csr_readdata),                      //  output,   width = 32,                               .readdata
		.pb_mm_bridge_address                     (pb_mm_bridge_address),                                                   //   input,   width = 17,                   pb_mm_bridge.address
		.pb_mm_bridge_chipselect                  (pb_mm_bridge_chipselect),                                                //   input,    width = 1,                               .chipselect
		.pb_mm_bridge_read                        (pb_mm_bridge_read),                                                      //   input,    width = 1,                               .read
		.pb_mm_bridge_readdata                    (pb_mm_bridge_readdata),                                                  //  output,   width = 32,                               .readdata
		.pb_mm_bridge_write                       (pb_mm_bridge_write),                                                     //   input,    width = 1,                               .write
		.pb_mm_bridge_writedata                   (pb_mm_bridge_writedata),                                                 //   input,   width = 32,                               .writedata
		.pb_mm_bridge_byteenable                  (pb_mm_bridge_byteenable),                                                //   input,    width = 4,                               .byteenable
		.pb_mm_bridge_waitrequest                 (pb_mm_bridge_waitrequest),                                               //  output,    width = 1,                               .waitrequest
		.lphy_ss_config_csr_address               (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_address),               //   input,    width = 8,             lphy_ss_config_csr.address
		.lphy_ss_config_csr_write                 (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_write),                 //   input,    width = 1,                               .write
		.lphy_ss_config_csr_writedata             (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_writedata),             //   input,   width = 32,                               .writedata
		.lphy_ss_config_csr_readdata              (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_readdata),              //  output,   width = 32,                               .readdata
		.lphy_ss_config_csr_read                  (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_read),                  //   input,    width = 1,                               .read
		.lphy_ss_config_csr_waitrequest           (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_waitrequest),           //  output,    width = 1,                               .waitrequest
		.lphy_ss_config_csr_readdatavalid         (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_readdatavalid),         //  output,    width = 1,                               .readdatavalid
		.long_prach_lw_bridge_address_l2          (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_address),          //   input,    width = 4,        long_prach_lw_bridge_l2.address
		.long_prach_lw_bridge_write_l2            (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_write),            //   input,    width = 1,                               .write
		.long_prach_lw_bridge_readdata_l2         (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_readdata),         //  output,   width = 32,                               .readdata
		.long_prach_lw_bridge_writedata_l2        (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_writedata),        //   input,   width = 32,                               .writedata
		.long_prach_lw_bridge_waitrequest_l2      (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_waitrequest),      //  output,    width = 1,                               .waitrequest
		.long_prach_lw_bridge_readdatavalid_l2    (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_readdatavalid),    //  output,    width = 1,                               .readdatavalid
		.long_prach_lw_bridge_read_l2             (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_read),             //   input,    width = 1,                               .read
		.long_prach_lw_bridge_address_l1          (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_address),          //   input,    width = 4,        long_prach_lw_bridge_l1.address
		.long_prach_lw_bridge_write_l1            (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_write),            //   input,    width = 1,                               .write
		.long_prach_lw_bridge_readdata_l1         (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_readdata),         //  output,   width = 32,                               .readdata
		.long_prach_lw_bridge_writedata_l1        (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_writedata),        //   input,   width = 32,                               .writedata
		.long_prach_lw_bridge_waitrequest_l1      (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_waitrequest),      //  output,    width = 1,                               .waitrequest
		.long_prach_lw_bridge_readdatavalid_l1    (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_readdatavalid),    //  output,    width = 1,                               .readdatavalid
		.long_prach_lw_bridge_read_l1             (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_read),             //   input,    width = 1,                               .read
		.short_prach2_busIn_writedata             (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_writedata),       //   input,   width = 32,       short_prach_lw_bridge_l2.writedata
		.short_prach2_busIn_address               (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_address),         //   input,   width = 10,                               .address
		.short_prach2_busIn_write                 (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_write),           //   input,    width = 1,                               .write
		.short_prach2_busIn_read                  (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_read),            //   input,    width = 1,                               .read
		.short_prach2_busOut_readdatavalid        (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_readdatavalid),   //  output,    width = 1,                               .readdatavalid
		.short_prach2_busOut_readdata             (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_readdata),        //  output,   width = 32,                               .readdata
		.short_prach2_busOut_waitrequest          (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_waitrequest),     //  output,    width = 1,                               .waitrequest
		.short_prach1_busIn_writedata             (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_writedata),       //   input,   width = 32,       short_prach_lw_bridge_l1.writedata
		.short_prach1_busIn_address               (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_address),         //   input,   width = 10,                               .address
		.short_prach1_busIn_write                 (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_write),           //   input,    width = 1,                               .write
		.short_prach1_busIn_read                  (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_read),            //   input,    width = 1,                               .read
		.short_prach1_busOut_readdatavalid        (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_readdatavalid),   //  output,    width = 1,                               .readdatavalid
		.short_prach1_busOut_readdata             (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_readdata),        //  output,   width = 32,                               .readdata
		.short_prach1_busOut_waitrequest          (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_waitrequest),     //  output,    width = 1,                               .waitrequest
		.clk_dsp                                  (clk_dsp_out_clk_clk),                                                    //   input,    width = 1,                      clock_dsp.clk
		.clk_csr                                  (clk_csr_out_clk_clk),                                                    //   input,    width = 1,                      clock_csr.clk
		.clk_eth_xran_dl                          (clk_xran_dl_out_clk_clk),                                                //   input,    width = 1,              clock_eth_xran_dl.clk
		.clk_eth_xran_ul                          (clk_xran_ul_out_clk_clk),                                                //   input,    width = 1,              clock_eth_xran_ul.clk
		.rst_dsp_n                                (reset_dsp_out_reset_reset),                                              //   input,    width = 1,                    reset_dsp_n.reset_n
		.rst_csr_n                                (~reset_csr_out_reset_reset),                                             //   input,    width = 1,                    reset_csr_n.reset_n
		.rst_eth_xran_n_dl                        (reset_xran_dl_out_reset_reset),                                          //   input,    width = 1,            reset_eth_xran_dl_n.reset_n
		.rst_eth_xran_n_ul                        (reset_xran_ul_out_reset_reset),                                          //   input,    width = 1,            reset_eth_xran_ul_n.reset_n
		.xran_demapper_source_valid               (xran_demapper_source_valid),                                             //   input,    width = 1,           xran_demapper_source.valid
		.xran_demapper_source_data                (xran_demapper_source_data),                                              //   input,  width = 128,                               .data
		.xran_demapper_source_endofpacket         (xran_demapper_source_endofpacket),                                       //   input,    width = 1,                               .endofpacket
		.xran_demapper_source_startofpacket       (xran_demapper_source_startofpacket),                                     //   input,    width = 1,                               .startofpacket
		.xran_demapper_source_ready               (xran_demapper_source_ready),                                             //  output,    width = 1,                               .ready
		.xran_demapper_source_channel             (xran_demapper_source_channel),                                           //   input,   width = 16,                               .channel
		.ifft_source_valid1                       (ifft_source_l1_valid),                                                   //  output,    width = 1,                 ifft_source_l1.valid
		.ifft_source_data1                        (ifft_source_l1_data),                                                    //  output,   width = 32,                               .data
		.ifft_source_channel1                     (ifft_source_l1_channel),                                                 //  output,    width = 8,                               .channel
		.ifft_source_valid2                       (ifft_source_l2_valid),                                                   //  output,    width = 1,                 ifft_source_l2.valid
		.ifft_source_data2                        (ifft_source_l2_data),                                                    //  output,   width = 32,                               .data
		.ifft_source_channel2                     (ifft_source_l2_channel),                                                 //  output,    width = 8,                               .channel
		.coupling_pusch_avst_sink_valid_l1        (coupling_pusch_avst_sink_l1_valid),                                      //  output,    width = 1,    coupling_pusch_avst_sink_l1.valid
		.coupling_pusch_avst_sink_data_l1         (coupling_pusch_avst_sink_l1_data),                                       //  output,   width = 32,                               .data
		.coupling_pusch_avst_sink_channel_l1      (coupling_pusch_avst_sink_l1_channel),                                    //  output,   width = 16,                               .channel
		.coupling_pusch_avst_sink_sop_l1          (coupling_pusch_avst_sink_l1_startofpacket),                              //  output,    width = 1,                               .startofpacket
		.coupling_pusch_avst_sink_eop_l1          (coupling_pusch_avst_sink_l1_endofpacket),                                //  output,    width = 1,                               .endofpacket
		.coupling_pusch_avst_sink_valid_l2        (coupling_pusch_avst_sink_l2_valid),                                      //  output,    width = 1,    coupling_pusch_avst_sink_l2.valid
		.coupling_pusch_avst_sink_data_l2         (coupling_pusch_avst_sink_l2_data),                                       //  output,   width = 32,                               .data
		.coupling_pusch_avst_sink_channel_l2      (coupling_pusch_avst_sink_l2_channel),                                    //  output,   width = 16,                               .channel
		.coupling_pusch_avst_sink_sop_l2          (coupling_pusch_avst_sink_l2_startofpacket),                              //  output,    width = 1,                               .startofpacket
		.coupling_pusch_avst_sink_eop_l2          (coupling_pusch_avst_sink_l2_endofpacket),                                //  output,    width = 1,                               .endofpacket
		.coupling_prach_avst_sink_valid_l1        (coupling_prach_avst_sink_l1_valid),                                      //  output,    width = 1,    coupling_prach_avst_sink_l1.valid
		.coupling_prach_avst_sink_data_l1         (coupling_prach_avst_sink_l1_data),                                       //  output,   width = 32,                               .data
		.coupling_prach_avst_sink_channel_l1      (coupling_prach_avst_sink_l1_channel),                                    //  output,   width = 16,                               .channel
		.coupling_prach_avst_sink_sop_l1          (coupling_prach_avst_sink_l1_startofpacket),                              //  output,    width = 1,                               .startofpacket
		.coupling_prach_avst_sink_eop_l1          (coupling_prach_avst_sink_l1_endofpacket),                                //  output,    width = 1,                               .endofpacket
		.coupling_prach_avst_sink_valid_l2        (coupling_prach_avst_sink_l2_valid),                                      //  output,    width = 1,    coupling_prach_avst_sink_l2.valid
		.coupling_prach_avst_sink_data_l2         (coupling_prach_avst_sink_l2_data),                                       //  output,   width = 32,                               .data
		.coupling_prach_avst_sink_channel_l2      (coupling_prach_avst_sink_l2_channel),                                    //  output,   width = 16,                               .channel
		.coupling_prach_avst_sink_sop_l2          (coupling_prach_avst_sink_l2_startofpacket),                              //  output,    width = 1,                               .startofpacket
		.coupling_prach_avst_sink_eop_l2          (coupling_prach_avst_sink_l2_endofpacket),                                //  output,    width = 1,                               .endofpacket
		.xran_demapper_cplane_valid               (xran_demapper_cplane_source_valid),                                      //   input,    width = 1,    xran_demapper_cplane_source.valid
		.xran_demapper_cplane_startofpacket       (xran_demapper_cplane_source_startofpacket),                              //   input,    width = 1,                               .startofpacket
		.xran_demapper_cplane_endofpacket         (xran_demapper_cplane_source_endofpacket),                                //   input,    width = 1,                               .endofpacket
		.pb_avst_sink_valid                       (pb_avst_sink_valid),                                                     //   input,    width = 1,                   pb_avst_sink.valid
		.pb_avst_sink_data                        (pb_avst_sink_data),                                                      //   input,   width = 64,                               .data
		.pb_avst_sink_ready                       (pb_avst_sink_ready),                                                     //  output,    width = 1,                               .ready
		.bw_config_cc1                            (bw_confg_cc1_bw_config_cc1),                                             //  output,    width = 8,                   bw_confg_cc1.bw_config_cc1
		.bw_config_cc2                            (bw_confg_cc2_bw_config_cc2),                                             //  output,    width = 8,                   bw_confg_cc2.bw_config_cc2
		.radio_config_status                      (radio_config_status_radio_config_status),                                //  output,   width = 56,            radio_config_status.radio_config_status
		.short_long_prach_select                  (short_long_prach_select_data),                                           //  output,    width = 1,        short_long_prach_select.data
		.rx_rtc_id                                (rx_rtc_id_rx_rtc_id),                                                    //   input,   width = 16,                      rx_rtc_id.rx_rtc_id
		.rx_u_axc_id                              (rx_u_axc_id_rx_u_axc_id),                                                //   input,   width = 16,                    rx_u_axc_id.rx_u_axc_id
		.rx_rtc_id_dl                             (rx_rtc_id_dl_rx_rtc_id_dl),                                              //   input,   width = 16,                   rx_rtc_id_dl.rx_rtc_id_dl
		.lphy_ss_ul_sink_valid1                   (lphy_ss_ul_sink_l1_valid),                                               //   input,    width = 1,             lphy_ss_ul_sink_l1.valid
		.lphy_ss_ul_sink_data1                    (lphy_ss_ul_sink_l1_data),                                                //   input,   width = 32,                               .data
		.lphy_ss_ul_sink_channel1                 (lphy_ss_ul_sink_l1_channel),                                             //   input,    width = 8,                               .channel
		.lphy_ss_ul_sink_valid2                   (lphy_ss_ul_sink_l2_valid),                                               //   input,    width = 1,             lphy_ss_ul_sink_l2.valid
		.lphy_ss_ul_sink_data2                    (lphy_ss_ul_sink_l2_data),                                                //   input,   width = 32,                               .data
		.lphy_ss_ul_sink_channel2                 (lphy_ss_ul_sink_l2_channel),                                             //   input,    width = 8,                               .channel
		.rst_soft_n                               (rst_soft_n_rst_soft_n),                                                  //  output,    width = 1,                     rst_soft_n.rst_soft_n
		.coupling_pusch_timing_ref                (coupling_pusch_timing_ref_data),                                         //  output,   width = 32,      coupling_pusch_timing_ref.data
		.coupling_prach_timing_ref                (coupling_prach_timing_ref_data),                                         //  output,   width = 32,      coupling_prach_timing_ref.data
		.oran_rx_cplane_concat                    (oran_rx_cplane_concat_data),                                             //   input,  width = 190,          oran_rx_cplane_concat.data
		.oran_rx_uplane_concat                    (oran_rx_uplane_concat_data),                                             //   input,   width = 68,          oran_rx_uplane_concat.data
		.lphy_avst_selctd_cap_intf_valid          (lphy_avst_selctd_cap_intf_valid),                                        //  output,    width = 1,      lphy_avst_selctd_cap_intf.valid
		.lphy_avst_selctd_cap_intf_data           (lphy_avst_selctd_cap_intf_data),                                         //  output,   width = 32,                               .data
		.lphy_avst_selctd_cap_intf_chan           (lphy_avst_selctd_cap_intf_channel),                                      //  output,    width = 3,                               .channel
		.ul_start_pulse_latch                     (ul_start_pulse_latch_data),                                              //  output,    width = 1,           ul_start_pulse_latch.data
		.frame_status_counter_reset               (frame_status_counter_reset_data),                                        //   input,    width = 1,     frame_status_counter_reset.data
		.interface_sel                            (lphy_ss_top_interface_sel_data),                                         //   input,   width = 32,                  interface_sel.data
		.dl_input_hfn_pulse                       (lphy_ss_top_dl_input_hfn_pulse_data),                                    //  output,    width = 1,             dl_input_hfn_pulse.data
		.pm_ifft_threash_mm_bridge_address_l1     (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_address),     //   input,    width = 6,   pm_ifft_threash_mm_bridge_l1.address
		.pm_ifft_threash_mm_bridge_chipselect_l1  (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_chipselect),  //   input,    width = 1,                               .chipselect
		.pm_ifft_threash_mm_bridge_read_l1        (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_read),        //   input,    width = 1,                               .read
		.pm_ifft_threash_mm_bridge_write_l1       (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_write),       //   input,    width = 1,                               .write
		.pm_ifft_threash_mm_bridge_writedata_l1   (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_writedata),   //   input,   width = 32,                               .writedata
		.pm_ifft_threash_mm_bridge_byteenable_l1  (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_byteenable),  //   input,    width = 4,                               .byteenable
		.pm_ifft_threash_mm_bridge_readdata_l1    (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_readdata),    //  output,   width = 32,                               .readdata
		.pm_ifft_threash_mm_bridge_waitrequest_l1 (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_waitrequest), //  output,    width = 1,                               .waitrequest
		.pwr_mtr_ifft_hist_done_intr_l1           (lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l1_irq),                         //  output,    width = 1, pwr_mtr_ifft_hist_done_intr_l1.irq
		.pwr_mtr_ifft_hist_done_intr_l2           (lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l2_irq),                         //  output,    width = 1, pwr_mtr_ifft_hist_done_intr_l2.irq
		.pm_ifft_threash_mm_bridge_address_l2     (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_address),     //   input,    width = 6,   pm_ifft_threash_mm_bridge_l2.address
		.pm_ifft_threash_mm_bridge_chipselect_l2  (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_chipselect),  //   input,    width = 1,                               .chipselect
		.pm_ifft_threash_mm_bridge_read_l2        (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_read),        //   input,    width = 1,                               .read
		.pm_ifft_threash_mm_bridge_write_l2       (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_write),       //   input,    width = 1,                               .write
		.pm_ifft_threash_mm_bridge_writedata_l2   (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_writedata),   //   input,   width = 32,                               .writedata
		.pm_ifft_threash_mm_bridge_byteenable_l2  (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_byteenable),  //   input,    width = 4,                               .byteenable
		.pm_ifft_threash_mm_bridge_readdata_l2    (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_readdata),    //  output,   width = 32,                               .readdata
		.pm_ifft_threash_mm_bridge_waitrequest_l2 (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_waitrequest), //  output,    width = 1,                               .waitrequest
		.pwr_mtr_ifft_config_csr_writedata_l1     (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_writedata),     //   input,   width = 32,     pwr_mtr_ifft_config_csr_l1.writedata
		.pwr_mtr_ifft_config_csr_read_l1          (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_read),          //   input,    width = 1,                               .read
		.pwr_mtr_ifft_config_csr_write_l1         (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_write),         //   input,    width = 1,                               .write
		.pwr_mtr_ifft_config_csr_readdata_l1      (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdata),      //  output,   width = 32,                               .readdata
		.pwr_mtr_ifft_config_csr_readdatavalid_l1 (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdatavalid), //  output,    width = 1,                               .readdatavalid
		.pwr_mtr_ifft_config_csr_address_l1       (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_address),       //   input,    width = 4,                               .address
		.pwr_mtr_ifft_config_csr_waitrequest_l1   (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_waitrequest),   //  output,    width = 1,                               .waitrequest
		.pwr_mtr_ifft_config_csr_writedata_l2     (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_writedata),     //   input,   width = 32,     pwr_mtr_ifft_config_csr_l2.writedata
		.pwr_mtr_ifft_config_csr_read_l2          (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_read),          //   input,    width = 1,                               .read
		.pwr_mtr_ifft_config_csr_write_l2         (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_write),         //   input,    width = 1,                               .write
		.pwr_mtr_ifft_config_csr_readdata_l2      (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdata),      //  output,   width = 32,                               .readdata
		.pwr_mtr_ifft_config_csr_readdatavalid_l2 (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdatavalid), //  output,    width = 1,                               .readdatavalid
		.pwr_mtr_ifft_config_csr_address_l2       (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_address),       //   input,    width = 4,                               .address
		.pwr_mtr_ifft_config_csr_waitrequest_l2   (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_waitrequest),   //  output,    width = 1,                               .waitrequest
		.pm_ifft_hist_mm_bridge_address_l1        (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_address),        //   input,   width = 12,      pm_ifft_hist_mm_bridge_l1.address
		.pm_ifft_hist_mm_bridge_chipselect_l1     (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_chipselect),     //   input,    width = 1,                               .chipselect
		.pm_ifft_hist_mm_bridge_read_l1           (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_read),           //   input,    width = 1,                               .read
		.pm_ifft_hist_mm_bridge_write_l1          (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_write),          //   input,    width = 1,                               .write
		.pm_ifft_hist_mm_bridge_writedata_l1      (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_writedata),      //   input,   width = 32,                               .writedata
		.pm_ifft_hist_mm_bridge_byteenable_l1     (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_byteenable),     //   input,    width = 4,                               .byteenable
		.pm_ifft_hist_mm_bridge_readdata_l1       (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdata),       //  output,   width = 32,                               .readdata
		.pm_ifft_hist_mm_bridge_readdatavalid_l1  (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdatavalid),  //  output,    width = 1,                               .readdatavalid
		.pm_ifft_hist_mm_bridge_waitrequest_l1    (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_waitrequest),    //  output,    width = 1,                               .waitrequest
		.pm_ifft_hist_mm_bridge_address_l2        (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_address),        //   input,   width = 12,      pm_ifft_hist_mm_bridge_l2.address
		.pm_ifft_hist_mm_bridge_chipselect_l2     (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_chipselect),     //   input,    width = 1,                               .chipselect
		.pm_ifft_hist_mm_bridge_read_l2           (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_read),           //   input,    width = 1,                               .read
		.pm_ifft_hist_mm_bridge_write_l2          (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_write),          //   input,    width = 1,                               .write
		.pm_ifft_hist_mm_bridge_writedata_l2      (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_writedata),      //   input,   width = 32,                               .writedata
		.pm_ifft_hist_mm_bridge_byteenable_l2     (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_byteenable),     //   input,    width = 4,                               .byteenable
		.pm_ifft_hist_mm_bridge_readdata_l2       (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdata),       //  output,   width = 32,                               .readdata
		.pm_ifft_hist_mm_bridge_readdatavalid_l2  (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdatavalid),  //  output,    width = 1,                               .readdatavalid
		.pm_ifft_hist_mm_bridge_waitrequest_l2    (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_waitrequest),    //  output,    width = 1,                               .waitrequest
		.pwr_mtr_fft_hist_done_intr_l1            (lphy_ss_top_pwr_mtr_fft_hist_done_intr_l1_irq),                          //  output,    width = 1,  pwr_mtr_fft_hist_done_intr_l1.irq
		.pwr_mtr_fft_hist_done_intr_l2            (lphy_ss_top_pwr_mtr_fft_hist_done_intr_l2_irq),                          //  output,    width = 1,  pwr_mtr_fft_hist_done_intr_l2.irq
		.duc_ddc_lpbk_en                          (lphy_ss_top_duc_ddc_lpbk_en_data),                                       //  output,    width = 1,                duc_ddc_lpbk_en.data
		.pm_fft_threash_mm_bridge_address_l1      (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_address),      //   input,    width = 6,    pm_fft_threash_mm_bridge_l1.address
		.pm_fft_threash_mm_bridge_chipselect_l1   (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_chipselect),   //   input,    width = 1,                               .chipselect
		.pm_fft_threash_mm_bridge_read_l1         (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_read),         //   input,    width = 1,                               .read
		.pm_fft_threash_mm_bridge_write_l1        (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_write),        //   input,    width = 1,                               .write
		.pm_fft_threash_mm_bridge_writedata_l1    (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_writedata),    //   input,   width = 32,                               .writedata
		.pm_fft_threash_mm_bridge_byteenable_l1   (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_byteenable),   //   input,    width = 4,                               .byteenable
		.pm_fft_threash_mm_bridge_readdata_l1     (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_readdata),     //  output,   width = 32,                               .readdata
		.pm_fft_threash_mm_bridge_waitrequest_l1  (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_waitrequest),  //  output,    width = 1,                               .waitrequest
		.pm_fft_threash_mm_bridge_address_l2      (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_address),      //   input,    width = 6,    pm_fft_threash_mm_bridge_l2.address
		.pm_fft_threash_mm_bridge_chipselect_l2   (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_chipselect),   //   input,    width = 1,                               .chipselect
		.pm_fft_threash_mm_bridge_read_l2         (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_read),         //   input,    width = 1,                               .read
		.pm_fft_threash_mm_bridge_write_l2        (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_write),        //   input,    width = 1,                               .write
		.pm_fft_threash_mm_bridge_writedata_l2    (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_writedata),    //   input,   width = 32,                               .writedata
		.pm_fft_threash_mm_bridge_byteenable_l2   (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_byteenable),   //   input,    width = 4,                               .byteenable
		.pm_fft_threash_mm_bridge_readdata_l2     (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_readdata),     //  output,   width = 32,                               .readdata
		.pm_fft_threash_mm_bridge_waitrequest_l2  (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_waitrequest),  //  output,    width = 1,                               .waitrequest
		.pwr_mtr_fft_config_csr_writedata_l1      (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_writedata),      //   input,   width = 32,      pwr_mtr_fft_config_csr_l1.writedata
		.pwr_mtr_fft_config_csr_read_l1           (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_read),           //   input,    width = 1,                               .read
		.pwr_mtr_fft_config_csr_write_l1          (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_write),          //   input,    width = 1,                               .write
		.pwr_mtr_fft_config_csr_readdata_l1       (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdata),       //  output,   width = 32,                               .readdata
		.pwr_mtr_fft_config_csr_readdatavalid_l1  (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdatavalid),  //  output,    width = 1,                               .readdatavalid
		.pwr_mtr_fft_config_csr_address_l1        (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_address),        //   input,    width = 4,                               .address
		.pwr_mtr_fft_config_csr_waitrequest_l1    (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_waitrequest),    //  output,    width = 1,                               .waitrequest
		.pwr_mtr_fft_config_csr_writedata_l2      (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_writedata),      //   input,   width = 32,      pwr_mtr_fft_config_csr_l2.writedata
		.pwr_mtr_fft_config_csr_read_l2           (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_read),           //   input,    width = 1,                               .read
		.pwr_mtr_fft_config_csr_write_l2          (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_write),          //   input,    width = 1,                               .write
		.pwr_mtr_fft_config_csr_readdata_l2       (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdata),       //  output,   width = 32,                               .readdata
		.pwr_mtr_fft_config_csr_readdatavalid_l2  (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdatavalid),  //  output,    width = 1,                               .readdatavalid
		.pwr_mtr_fft_config_csr_address_l2        (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_address),        //   input,    width = 4,                               .address
		.pwr_mtr_fft_config_csr_waitrequest_l2    (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_waitrequest),    //  output,    width = 1,                               .waitrequest
		.pm_fft_hist_mm_bridge_address_l1         (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_address),         //   input,   width = 12,       pm_fft_hist_mm_bridge_l1.address
		.pm_fft_hist_mm_bridge_chipselect_l1      (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_chipselect),      //   input,    width = 1,                               .chipselect
		.pm_fft_hist_mm_bridge_read_l1            (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_read),            //   input,    width = 1,                               .read
		.pm_fft_hist_mm_bridge_write_l1           (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_write),           //   input,    width = 1,                               .write
		.pm_fft_hist_mm_bridge_writedata_l1       (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_writedata),       //   input,   width = 32,                               .writedata
		.pm_fft_hist_mm_bridge_byteenable_l1      (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_byteenable),      //   input,    width = 4,                               .byteenable
		.pm_fft_hist_mm_bridge_readdata_l1        (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdata),        //  output,   width = 32,                               .readdata
		.pm_fft_hist_mm_bridge_readdatavalid_l1   (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdatavalid),   //  output,    width = 1,                               .readdatavalid
		.pm_fft_hist_mm_bridge_waitrequest_l1     (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_waitrequest),     //  output,    width = 1,                               .waitrequest
		.pm_fft_hist_mm_bridge_address_l2         (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_address),         //   input,   width = 12,       pm_fft_hist_mm_bridge_l2.address
		.pm_fft_hist_mm_bridge_chipselect_l2      (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_chipselect),      //   input,    width = 1,                               .chipselect
		.pm_fft_hist_mm_bridge_read_l2            (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_read),            //   input,    width = 1,                               .read
		.pm_fft_hist_mm_bridge_write_l2           (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_write),           //   input,    width = 1,                               .write
		.pm_fft_hist_mm_bridge_writedata_l2       (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_writedata),       //   input,   width = 32,                               .writedata
		.pm_fft_hist_mm_bridge_byteenable_l2      (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_byteenable),      //   input,    width = 4,                               .byteenable
		.pm_fft_hist_mm_bridge_readdata_l2        (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdata),        //  output,   width = 32,                               .readdata
		.pm_fft_hist_mm_bridge_readdatavalid_l2   (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdatavalid),   //  output,    width = 1,                               .readdatavalid
		.pm_fft_hist_mm_bridge_waitrequest_l2     (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_waitrequest),     //  output,    width = 1,                               .waitrequest
		.pm_stat_ifft_mm_bridge_address_l1        (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_address),        //   input,   width = 10,      pm_stat_ifft_mm_bridge_l1.address
		.pm_stat_ifft_mm_bridge_chipselect_l1     (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_chipselect),     //   input,    width = 1,                               .chipselect
		.pm_stat_ifft_mm_bridge_read_l1           (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_read),           //   input,    width = 1,                               .read
		.pm_stat_ifft_mm_bridge_write_l1          (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_write),          //   input,    width = 1,                               .write
		.pm_stat_ifft_mm_bridge_writedata_l1      (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_writedata),      //   input,   width = 32,                               .writedata
		.pm_stat_ifft_mm_bridge_byteenable_l1     (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_byteenable),     //   input,    width = 4,                               .byteenable
		.pm_stat_ifft_mm_bridge_readdata_l1       (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdata),       //  output,   width = 32,                               .readdata
		.pm_stat_ifft_mm_bridge_readdatavalid_l1  (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdatavalid),  //  output,    width = 1,                               .readdatavalid
		.pm_stat_ifft_mm_bridge_waitrequest_l1    (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_waitrequest),    //  output,    width = 1,                               .waitrequest
		.pm_stat_ifft_mm_bridge_address_l2        (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_address),        //   input,   width = 10,      pm_stat_ifft_mm_bridge_l2.address
		.pm_stat_ifft_mm_bridge_chipselect_l2     (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_chipselect),     //   input,    width = 1,                               .chipselect
		.pm_stat_ifft_mm_bridge_read_l2           (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_read),           //   input,    width = 1,                               .read
		.pm_stat_ifft_mm_bridge_write_l2          (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_write),          //   input,    width = 1,                               .write
		.pm_stat_ifft_mm_bridge_writedata_l2      (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_writedata),      //   input,   width = 32,                               .writedata
		.pm_stat_ifft_mm_bridge_byteenable_l2     (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_byteenable),     //   input,    width = 4,                               .byteenable
		.pm_stat_ifft_mm_bridge_readdata_l2       (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdata),       //  output,   width = 32,                               .readdata
		.pm_stat_ifft_mm_bridge_readdatavalid_l2  (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdatavalid),  //  output,    width = 1,                               .readdatavalid
		.pm_stat_ifft_mm_bridge_waitrequest_l2    (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_waitrequest),    //  output,    width = 1,                               .waitrequest
		.pm_stat_fft_mm_bridge_address_l1         (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_address),         //   input,   width = 10,       pm_stat_fft_mm_bridge_l1.address
		.pm_stat_fft_mm_bridge_chipselect_l1      (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_chipselect),      //   input,    width = 1,                               .chipselect
		.pm_stat_fft_mm_bridge_read_l1            (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_read),            //   input,    width = 1,                               .read
		.pm_stat_fft_mm_bridge_write_l1           (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_write),           //   input,    width = 1,                               .write
		.pm_stat_fft_mm_bridge_writedata_l1       (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_writedata),       //   input,   width = 32,                               .writedata
		.pm_stat_fft_mm_bridge_byteenable_l1      (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_byteenable),      //   input,    width = 4,                               .byteenable
		.pm_stat_fft_mm_bridge_readdata_l1        (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdata),        //  output,   width = 32,                               .readdata
		.pm_stat_fft_mm_bridge_readdatavalid_l1   (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdatavalid),   //  output,    width = 1,                               .readdatavalid
		.pm_stat_fft_mm_bridge_waitrequest_l1     (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_waitrequest),     //  output,    width = 1,                               .waitrequest
		.pm_stat_fft_mm_bridge_address_l2         (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_address),         //   input,   width = 10,       pm_stat_fft_mm_bridge_l2.address
		.pm_stat_fft_mm_bridge_chipselect_l2      (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_chipselect),      //   input,    width = 1,                               .chipselect
		.pm_stat_fft_mm_bridge_read_l2            (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_read),            //   input,    width = 1,                               .read
		.pm_stat_fft_mm_bridge_write_l2           (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_write),           //   input,    width = 1,                               .write
		.pm_stat_fft_mm_bridge_writedata_l2       (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_writedata),       //   input,   width = 32,                               .writedata
		.pm_stat_fft_mm_bridge_byteenable_l2      (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_byteenable),      //   input,    width = 4,                               .byteenable
		.pm_stat_fft_mm_bridge_readdata_l2        (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdata),        //  output,   width = 32,                               .readdata
		.pm_stat_fft_mm_bridge_readdatavalid_l2   (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdatavalid),   //  output,    width = 1,                               .readdatavalid
		.pm_stat_fft_mm_bridge_waitrequest_l2     (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_waitrequest)      //  output,    width = 1,                               .waitrequest
	);

	lphy_ss_reset_csr reset_csr (
		.clk       (clk_csr_out_clk_clk),       //   input,  width = 1,       clk.clk
		.in_reset  (reset_csr_reset),           //   input,  width = 1,  in_reset.reset
		.out_reset (reset_csr_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	lphy_ss_reset_dsp reset_dsp (
		.clk         (clk_dsp_out_clk_clk),       //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_dsp_in_reset_n),      //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (reset_dsp_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	lphy_ss_reset_xran_dl reset_xran_dl (
		.clk         (clk_xran_dl_out_clk_clk),       //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_xran_dl_reset_n),         //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (reset_xran_dl_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	lphy_ss_reset_xran_ul reset_xran_ul (
		.clk         (clk_xran_ul_out_clk_clk),       //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_xran_ul_reset_n),         //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (reset_xran_ul_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	lphy_ss_top_altera_mm_interconnect_1920_zqsa5uq mm_interconnect_0 (
		.h2f_lw_bridge_m0_address                                      (h2f_lw_bridge_m0_address),                                               //   input,  width = 19,                                        h2f_lw_bridge_m0.address
		.h2f_lw_bridge_m0_waitrequest                                  (h2f_lw_bridge_m0_waitrequest),                                           //  output,   width = 1,                                                        .waitrequest
		.h2f_lw_bridge_m0_burstcount                                   (h2f_lw_bridge_m0_burstcount),                                            //   input,   width = 1,                                                        .burstcount
		.h2f_lw_bridge_m0_byteenable                                   (h2f_lw_bridge_m0_byteenable),                                            //   input,   width = 4,                                                        .byteenable
		.h2f_lw_bridge_m0_read                                         (h2f_lw_bridge_m0_read),                                                  //   input,   width = 1,                                                        .read
		.h2f_lw_bridge_m0_readdata                                     (h2f_lw_bridge_m0_readdata),                                              //  output,  width = 32,                                                        .readdata
		.h2f_lw_bridge_m0_readdatavalid                                (h2f_lw_bridge_m0_readdatavalid),                                         //  output,   width = 1,                                                        .readdatavalid
		.h2f_lw_bridge_m0_write                                        (h2f_lw_bridge_m0_write),                                                 //   input,   width = 1,                                                        .write
		.h2f_lw_bridge_m0_writedata                                    (h2f_lw_bridge_m0_writedata),                                             //   input,  width = 32,                                                        .writedata
		.h2f_lw_bridge_m0_debugaccess                                  (h2f_lw_bridge_m0_debugaccess),                                           //   input,   width = 1,                                                        .debugaccess
		.lphy_ss_top_fft1_busin_address                                (mm_interconnect_0_lphy_ss_top_fft1_busin_address),                       //  output,  width = 14,                                  lphy_ss_top_fft1_busin.address
		.lphy_ss_top_fft1_busin_write                                  (mm_interconnect_0_lphy_ss_top_fft1_busin_write),                         //  output,   width = 1,                                                        .write
		.lphy_ss_top_fft1_busin_read                                   (mm_interconnect_0_lphy_ss_top_fft1_busin_read),                          //  output,   width = 1,                                                        .read
		.lphy_ss_top_fft1_busin_readdata                               (mm_interconnect_0_lphy_ss_top_fft1_busin_readdata),                      //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_fft1_busin_writedata                              (mm_interconnect_0_lphy_ss_top_fft1_busin_writedata),                     //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_fft1_busin_readdatavalid                          (mm_interconnect_0_lphy_ss_top_fft1_busin_readdatavalid),                 //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_fft1_busin_waitrequest                            (mm_interconnect_0_lphy_ss_top_fft1_busin_waitrequest),                   //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_fft2_busin_address                                (mm_interconnect_0_lphy_ss_top_fft2_busin_address),                       //  output,  width = 14,                                  lphy_ss_top_fft2_busin.address
		.lphy_ss_top_fft2_busin_write                                  (mm_interconnect_0_lphy_ss_top_fft2_busin_write),                         //  output,   width = 1,                                                        .write
		.lphy_ss_top_fft2_busin_read                                   (mm_interconnect_0_lphy_ss_top_fft2_busin_read),                          //  output,   width = 1,                                                        .read
		.lphy_ss_top_fft2_busin_readdata                               (mm_interconnect_0_lphy_ss_top_fft2_busin_readdata),                      //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_fft2_busin_writedata                              (mm_interconnect_0_lphy_ss_top_fft2_busin_writedata),                     //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_fft2_busin_readdatavalid                          (mm_interconnect_0_lphy_ss_top_fft2_busin_readdatavalid),                 //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_fft2_busin_waitrequest                            (mm_interconnect_0_lphy_ss_top_fft2_busin_waitrequest),                   //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_ifft1_busin_address                               (mm_interconnect_0_lphy_ss_top_ifft1_busin_address),                      //  output,  width = 14,                                 lphy_ss_top_ifft1_busin.address
		.lphy_ss_top_ifft1_busin_write                                 (mm_interconnect_0_lphy_ss_top_ifft1_busin_write),                        //  output,   width = 1,                                                        .write
		.lphy_ss_top_ifft1_busin_read                                  (mm_interconnect_0_lphy_ss_top_ifft1_busin_read),                         //  output,   width = 1,                                                        .read
		.lphy_ss_top_ifft1_busin_readdata                              (mm_interconnect_0_lphy_ss_top_ifft1_busin_readdata),                     //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_ifft1_busin_writedata                             (mm_interconnect_0_lphy_ss_top_ifft1_busin_writedata),                    //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_ifft1_busin_readdatavalid                         (mm_interconnect_0_lphy_ss_top_ifft1_busin_readdatavalid),                //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_ifft1_busin_waitrequest                           (mm_interconnect_0_lphy_ss_top_ifft1_busin_waitrequest),                  //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_ifft2_busin_address                               (mm_interconnect_0_lphy_ss_top_ifft2_busin_address),                      //  output,  width = 14,                                 lphy_ss_top_ifft2_busin.address
		.lphy_ss_top_ifft2_busin_write                                 (mm_interconnect_0_lphy_ss_top_ifft2_busin_write),                        //  output,   width = 1,                                                        .write
		.lphy_ss_top_ifft2_busin_read                                  (mm_interconnect_0_lphy_ss_top_ifft2_busin_read),                         //  output,   width = 1,                                                        .read
		.lphy_ss_top_ifft2_busin_readdata                              (mm_interconnect_0_lphy_ss_top_ifft2_busin_readdata),                     //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_ifft2_busin_writedata                             (mm_interconnect_0_lphy_ss_top_ifft2_busin_writedata),                    //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_ifft2_busin_readdatavalid                         (mm_interconnect_0_lphy_ss_top_ifft2_busin_readdatavalid),                //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_ifft2_busin_waitrequest                           (mm_interconnect_0_lphy_ss_top_ifft2_busin_waitrequest),                  //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_long_prach_lw_bridge_l1_address                   (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_address),          //  output,   width = 4,                     lphy_ss_top_long_prach_lw_bridge_l1.address
		.lphy_ss_top_long_prach_lw_bridge_l1_write                     (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_write),            //  output,   width = 1,                                                        .write
		.lphy_ss_top_long_prach_lw_bridge_l1_read                      (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_read),             //  output,   width = 1,                                                        .read
		.lphy_ss_top_long_prach_lw_bridge_l1_readdata                  (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_readdata),         //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_long_prach_lw_bridge_l1_writedata                 (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_writedata),        //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_long_prach_lw_bridge_l1_readdatavalid             (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_readdatavalid),    //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_long_prach_lw_bridge_l1_waitrequest               (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l1_waitrequest),      //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_long_prach_lw_bridge_l2_address                   (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_address),          //  output,   width = 4,                     lphy_ss_top_long_prach_lw_bridge_l2.address
		.lphy_ss_top_long_prach_lw_bridge_l2_write                     (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_write),            //  output,   width = 1,                                                        .write
		.lphy_ss_top_long_prach_lw_bridge_l2_read                      (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_read),             //  output,   width = 1,                                                        .read
		.lphy_ss_top_long_prach_lw_bridge_l2_readdata                  (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_readdata),         //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_long_prach_lw_bridge_l2_writedata                 (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_writedata),        //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_long_prach_lw_bridge_l2_readdatavalid             (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_readdatavalid),    //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_long_prach_lw_bridge_l2_waitrequest               (mm_interconnect_0_lphy_ss_top_long_prach_lw_bridge_l2_waitrequest),      //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_lphy_ss_config_csr_address                        (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_address),               //  output,   width = 8,                          lphy_ss_top_lphy_ss_config_csr.address
		.lphy_ss_top_lphy_ss_config_csr_write                          (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_write),                 //  output,   width = 1,                                                        .write
		.lphy_ss_top_lphy_ss_config_csr_read                           (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_read),                  //  output,   width = 1,                                                        .read
		.lphy_ss_top_lphy_ss_config_csr_readdata                       (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_readdata),              //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_lphy_ss_config_csr_writedata                      (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_writedata),             //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_lphy_ss_config_csr_readdatavalid                  (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_readdatavalid),         //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_lphy_ss_config_csr_waitrequest                    (mm_interconnect_0_lphy_ss_top_lphy_ss_config_csr_waitrequest),           //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_pb_ddr_csr_address                                (mm_interconnect_0_lphy_ss_top_pb_ddr_csr_address),                       //  output,   width = 4,                                  lphy_ss_top_pb_ddr_csr.address
		.lphy_ss_top_pb_ddr_csr_write                                  (mm_interconnect_0_lphy_ss_top_pb_ddr_csr_write),                         //  output,   width = 1,                                                        .write
		.lphy_ss_top_pb_ddr_csr_readdata                               (mm_interconnect_0_lphy_ss_top_pb_ddr_csr_readdata),                      //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_pb_ddr_csr_writedata                              (mm_interconnect_0_lphy_ss_top_pb_ddr_csr_writedata),                     //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_pwr_mtr_fft_config_csr_l1_address                 (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_address),        //  output,   width = 4,                   lphy_ss_top_pwr_mtr_fft_config_csr_l1.address
		.lphy_ss_top_pwr_mtr_fft_config_csr_l1_write                   (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_write),          //  output,   width = 1,                                                        .write
		.lphy_ss_top_pwr_mtr_fft_config_csr_l1_read                    (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_read),           //  output,   width = 1,                                                        .read
		.lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdata                (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdata),       //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_pwr_mtr_fft_config_csr_l1_writedata               (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_writedata),      //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdatavalid           (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_readdatavalid),  //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_pwr_mtr_fft_config_csr_l1_waitrequest             (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l1_waitrequest),    //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_pwr_mtr_fft_config_csr_l2_address                 (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_address),        //  output,   width = 4,                   lphy_ss_top_pwr_mtr_fft_config_csr_l2.address
		.lphy_ss_top_pwr_mtr_fft_config_csr_l2_write                   (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_write),          //  output,   width = 1,                                                        .write
		.lphy_ss_top_pwr_mtr_fft_config_csr_l2_read                    (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_read),           //  output,   width = 1,                                                        .read
		.lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdata                (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdata),       //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_pwr_mtr_fft_config_csr_l2_writedata               (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_writedata),      //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdatavalid           (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_readdatavalid),  //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_pwr_mtr_fft_config_csr_l2_waitrequest             (mm_interconnect_0_lphy_ss_top_pwr_mtr_fft_config_csr_l2_waitrequest),    //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l1_address                (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_address),       //  output,   width = 4,                  lphy_ss_top_pwr_mtr_ifft_config_csr_l1.address
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l1_write                  (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_write),         //  output,   width = 1,                                                        .write
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l1_read                   (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_read),          //  output,   width = 1,                                                        .read
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdata               (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdata),      //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l1_writedata              (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_writedata),     //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdatavalid          (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_readdatavalid), //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l1_waitrequest            (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l1_waitrequest),   //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l2_address                (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_address),       //  output,   width = 4,                  lphy_ss_top_pwr_mtr_ifft_config_csr_l2.address
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l2_write                  (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_write),         //  output,   width = 1,                                                        .write
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l2_read                   (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_read),          //  output,   width = 1,                                                        .read
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdata               (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdata),      //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l2_writedata              (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_writedata),     //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdatavalid          (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_readdatavalid), //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_pwr_mtr_ifft_config_csr_l2_waitrequest            (mm_interconnect_0_lphy_ss_top_pwr_mtr_ifft_config_csr_l2_waitrequest),   //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_short_prach_lw_bridge_l1_address                  (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_address),         //  output,  width = 10,                    lphy_ss_top_short_prach_lw_bridge_l1.address
		.lphy_ss_top_short_prach_lw_bridge_l1_write                    (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_write),           //  output,   width = 1,                                                        .write
		.lphy_ss_top_short_prach_lw_bridge_l1_read                     (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_read),            //  output,   width = 1,                                                        .read
		.lphy_ss_top_short_prach_lw_bridge_l1_readdata                 (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_readdata),        //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_short_prach_lw_bridge_l1_writedata                (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_writedata),       //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_short_prach_lw_bridge_l1_readdatavalid            (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_readdatavalid),   //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_short_prach_lw_bridge_l1_waitrequest              (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l1_waitrequest),     //   input,   width = 1,                                                        .waitrequest
		.lphy_ss_top_short_prach_lw_bridge_l2_address                  (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_address),         //  output,  width = 10,                    lphy_ss_top_short_prach_lw_bridge_l2.address
		.lphy_ss_top_short_prach_lw_bridge_l2_write                    (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_write),           //  output,   width = 1,                                                        .write
		.lphy_ss_top_short_prach_lw_bridge_l2_read                     (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_read),            //  output,   width = 1,                                                        .read
		.lphy_ss_top_short_prach_lw_bridge_l2_readdata                 (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_readdata),        //   input,  width = 32,                                                        .readdata
		.lphy_ss_top_short_prach_lw_bridge_l2_writedata                (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_writedata),       //  output,  width = 32,                                                        .writedata
		.lphy_ss_top_short_prach_lw_bridge_l2_readdatavalid            (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_readdatavalid),   //   input,   width = 1,                                                        .readdatavalid
		.lphy_ss_top_short_prach_lw_bridge_l2_waitrequest              (mm_interconnect_0_lphy_ss_top_short_prach_lw_bridge_l2_waitrequest),     //   input,   width = 1,                                                        .waitrequest
		.h2f_lw_bridge_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                         //   input,   width = 1,               h2f_lw_bridge_reset_reset_bridge_in_reset.reset
		.h2f_lw_bridge_m0_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                         //   input,   width = 1, h2f_lw_bridge_m0_translator_reset_reset_bridge_in_reset.reset
		.clk_csr_out_clk_clk                                           (clk_csr_out_clk_clk)                                                     //   input,   width = 1,                                         clk_csr_out_clk.clk
	);

	lphy_ss_top_altera_mm_interconnect_1920_sjiabna mm_interconnect_1 (
		.h2f_bridge_m0_address                                      (h2f_bridge_m0_address),                                                  //   input,  width = 17,                                        h2f_bridge_m0.address
		.h2f_bridge_m0_waitrequest                                  (h2f_bridge_m0_waitrequest),                                              //  output,   width = 1,                                                     .waitrequest
		.h2f_bridge_m0_burstcount                                   (h2f_bridge_m0_burstcount),                                               //   input,   width = 1,                                                     .burstcount
		.h2f_bridge_m0_byteenable                                   (h2f_bridge_m0_byteenable),                                               //   input,   width = 4,                                                     .byteenable
		.h2f_bridge_m0_read                                         (h2f_bridge_m0_read),                                                     //   input,   width = 1,                                                     .read
		.h2f_bridge_m0_readdata                                     (h2f_bridge_m0_readdata),                                                 //  output,  width = 32,                                                     .readdata
		.h2f_bridge_m0_readdatavalid                                (h2f_bridge_m0_readdatavalid),                                            //  output,   width = 1,                                                     .readdatavalid
		.h2f_bridge_m0_write                                        (h2f_bridge_m0_write),                                                    //   input,   width = 1,                                                     .write
		.h2f_bridge_m0_writedata                                    (h2f_bridge_m0_writedata),                                                //   input,  width = 32,                                                     .writedata
		.h2f_bridge_m0_debugaccess                                  (h2f_bridge_m0_debugaccess),                                              //   input,   width = 1,                                                     .debugaccess
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_address               (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_address),         //  output,  width = 12,                 lphy_ss_top_pm_fft_hist_mm_bridge_l1.address
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_write                 (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_write),           //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_read                  (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_read),            //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdata              (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdata),        //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_writedata             (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_writedata),       //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_byteenable            (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_byteenable),      //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdatavalid         (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_readdatavalid),   //   input,   width = 1,                                                     .readdatavalid
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_waitrequest           (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_waitrequest),     //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_fft_hist_mm_bridge_l1_chipselect            (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l1_chipselect),      //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_address               (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_address),         //  output,  width = 12,                 lphy_ss_top_pm_fft_hist_mm_bridge_l2.address
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_write                 (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_write),           //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_read                  (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_read),            //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdata              (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdata),        //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_writedata             (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_writedata),       //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_byteenable            (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_byteenable),      //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdatavalid         (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_readdatavalid),   //   input,   width = 1,                                                     .readdatavalid
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_waitrequest           (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_waitrequest),     //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_fft_hist_mm_bridge_l2_chipselect            (mm_interconnect_1_lphy_ss_top_pm_fft_hist_mm_bridge_l2_chipselect),      //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_fft_threash_mm_bridge_l1_address            (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_address),      //  output,   width = 6,              lphy_ss_top_pm_fft_threash_mm_bridge_l1.address
		.lphy_ss_top_pm_fft_threash_mm_bridge_l1_write              (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_write),        //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_fft_threash_mm_bridge_l1_read               (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_read),         //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_fft_threash_mm_bridge_l1_readdata           (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_readdata),     //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_fft_threash_mm_bridge_l1_writedata          (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_writedata),    //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_fft_threash_mm_bridge_l1_byteenable         (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_byteenable),   //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_fft_threash_mm_bridge_l1_waitrequest        (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_waitrequest),  //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_fft_threash_mm_bridge_l1_chipselect         (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l1_chipselect),   //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_fft_threash_mm_bridge_l2_address            (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_address),      //  output,   width = 6,              lphy_ss_top_pm_fft_threash_mm_bridge_l2.address
		.lphy_ss_top_pm_fft_threash_mm_bridge_l2_write              (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_write),        //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_fft_threash_mm_bridge_l2_read               (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_read),         //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_fft_threash_mm_bridge_l2_readdata           (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_readdata),     //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_fft_threash_mm_bridge_l2_writedata          (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_writedata),    //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_fft_threash_mm_bridge_l2_byteenable         (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_byteenable),   //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_fft_threash_mm_bridge_l2_waitrequest        (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_waitrequest),  //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_fft_threash_mm_bridge_l2_chipselect         (mm_interconnect_1_lphy_ss_top_pm_fft_threash_mm_bridge_l2_chipselect),   //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_address              (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_address),        //  output,  width = 12,                lphy_ss_top_pm_ifft_hist_mm_bridge_l1.address
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_write                (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_write),          //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_read                 (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_read),           //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdata             (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdata),       //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_writedata            (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_writedata),      //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_byteenable           (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_byteenable),     //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdatavalid        (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_readdatavalid),  //   input,   width = 1,                                                     .readdatavalid
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_waitrequest          (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_waitrequest),    //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l1_chipselect           (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l1_chipselect),     //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_address              (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_address),        //  output,  width = 12,                lphy_ss_top_pm_ifft_hist_mm_bridge_l2.address
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_write                (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_write),          //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_read                 (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_read),           //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdata             (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdata),       //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_writedata            (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_writedata),      //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_byteenable           (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_byteenable),     //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdatavalid        (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_readdatavalid),  //   input,   width = 1,                                                     .readdatavalid
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_waitrequest          (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_waitrequest),    //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_ifft_hist_mm_bridge_l2_chipselect           (mm_interconnect_1_lphy_ss_top_pm_ifft_hist_mm_bridge_l2_chipselect),     //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l1_address           (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_address),     //  output,   width = 6,             lphy_ss_top_pm_ifft_threash_mm_bridge_l1.address
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l1_write             (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_write),       //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l1_read              (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_read),        //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l1_readdata          (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_readdata),    //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l1_writedata         (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_writedata),   //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l1_byteenable        (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_byteenable),  //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l1_waitrequest       (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_waitrequest), //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l1_chipselect        (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l1_chipselect),  //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l2_address           (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_address),     //  output,   width = 6,             lphy_ss_top_pm_ifft_threash_mm_bridge_l2.address
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l2_write             (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_write),       //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l2_read              (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_read),        //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l2_readdata          (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_readdata),    //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l2_writedata         (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_writedata),   //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l2_byteenable        (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_byteenable),  //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l2_waitrequest       (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_waitrequest), //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_ifft_threash_mm_bridge_l2_chipselect        (mm_interconnect_1_lphy_ss_top_pm_ifft_threash_mm_bridge_l2_chipselect),  //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_address               (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_address),         //  output,  width = 10,                 lphy_ss_top_pm_stat_fft_mm_bridge_l1.address
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_write                 (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_write),           //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_read                  (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_read),            //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdata              (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdata),        //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_writedata             (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_writedata),       //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_byteenable            (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_byteenable),      //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdatavalid         (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_readdatavalid),   //   input,   width = 1,                                                     .readdatavalid
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_waitrequest           (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_waitrequest),     //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_stat_fft_mm_bridge_l1_chipselect            (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l1_chipselect),      //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_address               (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_address),         //  output,  width = 10,                 lphy_ss_top_pm_stat_fft_mm_bridge_l2.address
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_write                 (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_write),           //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_read                  (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_read),            //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdata              (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdata),        //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_writedata             (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_writedata),       //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_byteenable            (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_byteenable),      //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdatavalid         (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_readdatavalid),   //   input,   width = 1,                                                     .readdatavalid
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_waitrequest           (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_waitrequest),     //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_stat_fft_mm_bridge_l2_chipselect            (mm_interconnect_1_lphy_ss_top_pm_stat_fft_mm_bridge_l2_chipselect),      //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_address              (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_address),        //  output,  width = 10,                lphy_ss_top_pm_stat_ifft_mm_bridge_l1.address
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_write                (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_write),          //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_read                 (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_read),           //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdata             (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdata),       //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_writedata            (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_writedata),      //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_byteenable           (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_byteenable),     //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdatavalid        (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_readdatavalid),  //   input,   width = 1,                                                     .readdatavalid
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_waitrequest          (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_waitrequest),    //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l1_chipselect           (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l1_chipselect),     //  output,   width = 1,                                                     .chipselect
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_address              (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_address),        //  output,  width = 10,                lphy_ss_top_pm_stat_ifft_mm_bridge_l2.address
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_write                (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_write),          //  output,   width = 1,                                                     .write
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_read                 (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_read),           //  output,   width = 1,                                                     .read
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdata             (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdata),       //   input,  width = 32,                                                     .readdata
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_writedata            (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_writedata),      //  output,  width = 32,                                                     .writedata
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_byteenable           (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_byteenable),     //  output,   width = 4,                                                     .byteenable
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdatavalid        (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_readdatavalid),  //   input,   width = 1,                                                     .readdatavalid
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_waitrequest          (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_waitrequest),    //   input,   width = 1,                                                     .waitrequest
		.lphy_ss_top_pm_stat_ifft_mm_bridge_l2_chipselect           (mm_interconnect_1_lphy_ss_top_pm_stat_ifft_mm_bridge_l2_chipselect),     //  output,   width = 1,                                                     .chipselect
		.h2f_bridge_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                         //   input,   width = 1,               h2f_bridge_reset_reset_bridge_in_reset.reset
		.h2f_bridge_m0_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                         //   input,   width = 1, h2f_bridge_m0_translator_reset_reset_bridge_in_reset.reset
		.clk_csr_out_clk_clk                                        (clk_csr_out_clk_clk)                                                     //   input,   width = 1,                                      clk_csr_out_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_csr_out_reset_reset),      //   input,  width = 1, reset_in0.reset
		.clk            (clk_csr_out_clk_clk),            //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

endmodule
