// qsys_top.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module qsys_top #(
		parameter FP_WIDTH = 32,
		parameter SIM_MODE = 0
	) (
		input  wire [19:0]  ftile_debug_status_econ_export,                                                          //                                                     ftile_debug_status_econ.export
		input  wire         hssi_ss_1_p0_axi_st_tx_reset_reset_n,                                                    //                                                hssi_ss_1_p0_axi_st_tx_reset.reset_n
		input  wire         hssi_ss_1_p0_axi_st_tx_interface_tvalid,                                                 //                                            hssi_ss_1_p0_axi_st_tx_interface.tvalid
		output wire         hssi_ss_1_p0_axi_st_tx_interface_tready,                                                 //                                                                            .tready
		input  wire [63:0]  hssi_ss_1_p0_axi_st_tx_interface_tdata,                                                  //                                                                            .tdata
		input  wire [7:0]   hssi_ss_1_p0_axi_st_tx_interface_tkeep,                                                  //                                                                            .tkeep
		input  wire         hssi_ss_1_p0_axi_st_tx_interface_tlast,                                                  //                                                                            .tlast
		input  wire [1:0]   hssi_ss_1_p0_axi_st_tx_interface_tuser,                                                  //                                                                            .tuser
		input  wire [93:0]  hssi_ss_1_p0_tx_tuser_ptp_tuser_1,                                                       //                                                   hssi_ss_1_p0_tx_tuser_ptp.tuser_1
		input  wire [327:0] hssi_ss_1_p0_tx_tuser_ptp_extended_tuser_2,                                              //                                          hssi_ss_1_p0_tx_tuser_ptp_extended.tuser_2
		input  wire         hssi_ss_1_p0_axi_st_tx_tuser_last_seg_interface_tx_last_segment,                         //                             hssi_ss_1_p0_axi_st_tx_tuser_last_seg_interface.tx_last_segment
		input  wire         hssi_ss_1_p0_axi_st_rx_reset_reset_n,                                                    //                                                hssi_ss_1_p0_axi_st_rx_reset.reset_n
		output wire [4:0]   hssi_ss_1_p0_rx_tuser_status_tuser_1,                                                    //                                                hssi_ss_1_p0_rx_tuser_status.tuser_1
		output wire         hssi_ss_1_p0_axi_st_tx_egrs0_interface_tvalid,                                           //                                      hssi_ss_1_p0_axi_st_tx_egrs0_interface.tvalid
		output wire [127:0] hssi_ss_1_p0_axi_st_tx_egrs0_interface_tdata,                                            //                                                                            .tdata
		output wire         hssi_ss_1_p0_axi_st_rx_ingrs0_interface_tvalid,                                          //                                     hssi_ss_1_p0_axi_st_rx_ingrs0_interface.tvalid
		output wire [95:0]  hssi_ss_1_p0_axi_st_rx_ingrs0_interface_tdata,                                           //                                                                            .tdata
		input  wire         hssi_ss_1_p0_tx_flow_control_interface_i_p0_tx_pause,                                    //                                      hssi_ss_1_p0_tx_flow_control_interface.i_p0_tx_pause
		input  wire [7:0]   hssi_ss_1_p0_tx_flow_control_interface_i_p0_tx_pfc,                                      //                                                                            .i_p0_tx_pfc
		output wire [0:0]   hssi_ss_1_p0_tx_srl_interface_p0_tx_serial,                                              //                                               hssi_ss_1_p0_tx_srl_interface.p0_tx_serial
		output wire [0:0]   hssi_ss_1_p0_tx_srl_interface_p0_tx_serial_n,                                            //                                                                            .p0_tx_serial_n
		input  wire [0:0]   hssi_ss_1_p0_rx_srl_interface_p0_rx_serial,                                              //                                               hssi_ss_1_p0_rx_srl_interface.p0_rx_serial
		input  wire [0:0]   hssi_ss_1_p0_rx_srl_interface_p0_rx_serial_n,                                            //                                                                            .p0_rx_serial_n
		output wire [2:0]   hssi_ss_1_p0_qsfp_led_sts_if_port0_led_speed,                                            //                                                hssi_ss_1_p0_qsfp_led_sts_if.port0_led_speed
		output wire [2:0]   hssi_ss_1_p0_qsfp_led_sts_if_port0_led_status,                                           //                                                                            .port0_led_status
		output wire [2:0]   hssi_ss_1_p1_qsfp_led_sts_if_port1_led_speed,                                            //                                                hssi_ss_1_p1_qsfp_led_sts_if.port1_led_speed
		output wire [2:0]   hssi_ss_1_p1_qsfp_led_sts_if_port1_led_status,                                           //                                                                            .port1_led_status
		output wire [2:0]   hssi_ss_1_p2_qsfp_led_sts_if_port2_led_speed,                                            //                                                hssi_ss_1_p2_qsfp_led_sts_if.port2_led_speed
		output wire [2:0]   hssi_ss_1_p2_qsfp_led_sts_if_port2_led_status,                                           //                                                                            .port2_led_status
		output wire [2:0]   hssi_ss_1_p3_qsfp_led_sts_if_port3_led_speed,                                            //                                                hssi_ss_1_p3_qsfp_led_sts_if.port3_led_speed
		output wire [2:0]   hssi_ss_1_p3_qsfp_led_sts_if_port3_led_status,                                           //                                                                            .port3_led_status
		output wire [2:0]   hssi_ss_1_p4_qsfp_led_sts_if_port4_led_speed,                                            //                                                hssi_ss_1_p4_qsfp_led_sts_if.port4_led_speed
		output wire [2:0]   hssi_ss_1_p4_qsfp_led_sts_if_port4_led_status,                                           //                                                                            .port4_led_status
		output wire [2:0]   hssi_ss_1_p5_qsfp_led_sts_if_port5_led_speed,                                            //                                                hssi_ss_1_p5_qsfp_led_sts_if.port5_led_speed
		output wire [2:0]   hssi_ss_1_p5_qsfp_led_sts_if_port5_led_status,                                           //                                                                            .port5_led_status
		output wire [2:0]   hssi_ss_1_p6_qsfp_led_sts_if_port6_led_speed,                                            //                                                hssi_ss_1_p6_qsfp_led_sts_if.port6_led_speed
		output wire [2:0]   hssi_ss_1_p6_qsfp_led_sts_if_port6_led_status,                                           //                                                                            .port6_led_status
		output wire [2:0]   hssi_ss_1_p7_qsfp_led_sts_if_port7_led_speed,                                            //                                                hssi_ss_1_p7_qsfp_led_sts_if.port7_led_speed
		output wire [2:0]   hssi_ss_1_p7_qsfp_led_sts_if_port7_led_status,                                           //                                                                            .port7_led_status
		output wire [2:0]   hssi_ss_1_p8_qsfp_led_sts_if_port8_led_speed,                                            //                                                hssi_ss_1_p8_qsfp_led_sts_if.port8_led_speed
		output wire [2:0]   hssi_ss_1_p8_qsfp_led_sts_if_port8_led_status,                                           //                                                                            .port8_led_status
		output wire [2:0]   hssi_ss_1_p9_qsfp_led_sts_if_port9_led_speed,                                            //                                                hssi_ss_1_p9_qsfp_led_sts_if.port9_led_speed
		output wire [2:0]   hssi_ss_1_p9_qsfp_led_sts_if_port9_led_status,                                           //                                                                            .port9_led_status
		output wire [2:0]   hssi_ss_1_p10_qsfp_led_sts_if_port10_led_speed,                                          //                                               hssi_ss_1_p10_qsfp_led_sts_if.port10_led_speed
		output wire [2:0]   hssi_ss_1_p10_qsfp_led_sts_if_port10_led_status,                                         //                                                                            .port10_led_status
		output wire [2:0]   hssi_ss_1_p11_qsfp_led_sts_if_port11_led_speed,                                          //                                               hssi_ss_1_p11_qsfp_led_sts_if.port11_led_speed
		output wire [2:0]   hssi_ss_1_p11_qsfp_led_sts_if_port11_led_status,                                         //                                                                            .port11_led_status
		output wire [2:0]   hssi_ss_1_p12_qsfp_led_sts_if_port12_led_speed,                                          //                                               hssi_ss_1_p12_qsfp_led_sts_if.port12_led_speed
		output wire [2:0]   hssi_ss_1_p12_qsfp_led_sts_if_port12_led_status,                                         //                                                                            .port12_led_status
		output wire [2:0]   hssi_ss_1_p13_qsfp_led_sts_if_port13_led_speed,                                          //                                               hssi_ss_1_p13_qsfp_led_sts_if.port13_led_speed
		output wire [2:0]   hssi_ss_1_p13_qsfp_led_sts_if_port13_led_status,                                         //                                                                            .port13_led_status
		output wire [2:0]   hssi_ss_1_p14_qsfp_led_sts_if_port14_led_speed,                                          //                                               hssi_ss_1_p14_qsfp_led_sts_if.port14_led_speed
		output wire [2:0]   hssi_ss_1_p14_qsfp_led_sts_if_port14_led_status,                                         //                                                                            .port14_led_status
		output wire [2:0]   hssi_ss_1_p15_qsfp_led_sts_if_port15_led_speed,                                          //                                               hssi_ss_1_p15_qsfp_led_sts_if.port15_led_speed
		output wire [2:0]   hssi_ss_1_p15_qsfp_led_sts_if_port15_led_status,                                         //                                                                            .port15_led_status
		output wire [2:0]   hssi_ss_1_p16_qsfp_led_sts_if_port16_led_speed,                                          //                                               hssi_ss_1_p16_qsfp_led_sts_if.port16_led_speed
		output wire [2:0]   hssi_ss_1_p16_qsfp_led_sts_if_port16_led_status,                                         //                                                                            .port16_led_status
		output wire [2:0]   hssi_ss_1_p17_qsfp_led_sts_if_port17_led_speed,                                          //                                               hssi_ss_1_p17_qsfp_led_sts_if.port17_led_speed
		output wire [2:0]   hssi_ss_1_p17_qsfp_led_sts_if_port17_led_status,                                         //                                                                            .port17_led_status
		output wire [2:0]   hssi_ss_1_p18_qsfp_led_sts_if_port18_led_speed,                                          //                                               hssi_ss_1_p18_qsfp_led_sts_if.port18_led_speed
		output wire [2:0]   hssi_ss_1_p18_qsfp_led_sts_if_port18_led_status,                                         //                                                                            .port18_led_status
		output wire [2:0]   hssi_ss_1_p19_qsfp_led_sts_if_port19_led_speed,                                          //                                               hssi_ss_1_p19_qsfp_led_sts_if.port19_led_speed
		output wire [2:0]   hssi_ss_1_p19_qsfp_led_sts_if_port19_led_status,                                         //                                                                            .port19_led_status
		output wire         hssi_ss_1_p0_misc_interface_p0_tx_lanes_stable,                                          //                                                 hssi_ss_1_p0_misc_interface.p0_tx_lanes_stable
		output wire         hssi_ss_1_p0_misc_interface_p0_rx_pcs_ready,                                             //                                                                            .p0_rx_pcs_ready
		output wire         hssi_ss_1_p0_misc_interface_o_p0_tx_pll_locked,                                          //                                                                            .o_p0_tx_pll_locked
		output wire         hssi_ss_1_p0_tx_ptp_ready_o_p0_tx_ptp_ready,                                             //                                                   hssi_ss_1_p0_tx_ptp_ready.o_p0_tx_ptp_ready
		output wire         hssi_ss_1_p0_rx_ptp_ready_o_p0_rx_ptp_ready,                                             //                                                   hssi_ss_1_p0_rx_ptp_ready.o_p0_rx_ptp_ready
		output wire         hssi_ss_1_p0_ptp_offset_data_valid_o_p0_rx_ptp_offset_data_valid,                        //                                          hssi_ss_1_p0_ptp_offset_data_valid.o_p0_rx_ptp_offset_data_valid
		output wire         hssi_ss_1_p0_ptp_offset_data_valid_o_p0_tx_ptp_offset_data_valid,                        //                                                                            .o_p0_tx_ptp_offset_data_valid
		input  wire         hssi_ss_1_subsystem_cold_rst_n_reset_n,                                                  //                                              hssi_ss_1_subsystem_cold_rst_n.reset_n
		output wire         hssi_ss_1_subsystem_cold_rst_ack_n_reset_n,                                              //                                          hssi_ss_1_subsystem_cold_rst_ack_n.reset_n
		input  wire         hssi_ss_1_i_p0_tx_rst_n_reset_n,                                                         //                                                     hssi_ss_1_i_p0_tx_rst_n.reset_n
		input  wire         hssi_ss_1_i_p0_rx_rst_n_reset_n,                                                         //                                                     hssi_ss_1_i_p0_rx_rst_n.reset_n
		output wire         hssi_ss_1_o_p0_rx_rst_ack_n_reset_n,                                                     //                                                 hssi_ss_1_o_p0_rx_rst_ack_n.reset_n
		output wire         hssi_ss_1_o_p0_tx_rst_ack_n_reset_n,                                                     //                                                 hssi_ss_1_o_p0_tx_rst_ack_n.reset_n
		input  wire [1:0]   hssi_ss_1_i_clk_ref_clk,                                                                 //                                                         hssi_ss_1_i_clk_ref.clk
		input  wire [1:0]   qsfpdd_status_pio_external_connection_export,                                            //                                       qsfpdd_status_pio_external_connection.export
		output wire [5:0]   qsfpdd_ctrl_pio_0_econ_export,                                                           //                                                      qsfpdd_ctrl_pio_0_econ.export
		input  wire         clk_csr_in_clk_clk,                                                                      //                                                              clk_csr_in_clk.clk
		input  wire         clk_dsp_in_clk_clk,                                                                      //                                                              clk_dsp_in_clk.clk
		output wire         hssi_ss_1_o_p0_clk_rec_div_clk,                                                          //                                                  hssi_ss_1_o_p0_clk_rec_div.clk
		output wire         ftile_out_clk_clk,                                                                       //                                                               ftile_out_clk.clk
		input  wire         dfd_subsystem_clock_bridge_dspby2_in_clk_clk,                                            //                                    dfd_subsystem_clock_bridge_dspby2_in_clk.clk
		input  wire         dma_subsys_ninit_done_reset,                                                             //                                                       dma_subsys_ninit_done.reset
		input  wire         dma_subsys_dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_valid,            //      dma_subsys_dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts.valid
		input  wire [95:0]  dma_subsys_dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_data,             //                                                                            .data
		input  wire [0:0]   ts_chs_compl_0_rst_bus_in_reset,                                                         //                                                   ts_chs_compl_0_rst_bus_in.reset
		input  wire [0:0]   dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_valid,            //      dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts.valid
		input  wire [19:0]  dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_fingerprint,      //                                                                            .fingerprint
		input  wire [95:0]  dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_data,             //                                                                            .data
		output wire         dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_valid,       // dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req.valid
		output wire [19:0]  dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_fingerprint, //                                                                            .fingerprint
		input  wire [43:0]  agilex_hps_f2h_stm_hw_events_stm_hwevents,                                               //                                                agilex_hps_f2h_stm_hw_events.stm_hwevents
		input  wire         agilex_hps_h2f_cs_ntrst,                                                                 //                                                           agilex_hps_h2f_cs.ntrst
		input  wire         agilex_hps_h2f_cs_tck,                                                                   //                                                                            .tck
		input  wire         agilex_hps_h2f_cs_tdi,                                                                   //                                                                            .tdi
		output wire         agilex_hps_h2f_cs_tdo,                                                                   //                                                                            .tdo
		output wire         agilex_hps_h2f_cs_tdoen,                                                                 //                                                                            .tdoen
		input  wire         agilex_hps_h2f_cs_tms,                                                                   //                                                                            .tms
		output wire         hps_io_EMAC1_TX_CLK,                                                                     //                                                                      hps_io.EMAC1_TX_CLK
		output wire         hps_io_EMAC1_TXD0,                                                                       //                                                                            .EMAC1_TXD0
		output wire         hps_io_EMAC1_TXD1,                                                                       //                                                                            .EMAC1_TXD1
		output wire         hps_io_EMAC1_TXD2,                                                                       //                                                                            .EMAC1_TXD2
		output wire         hps_io_EMAC1_TXD3,                                                                       //                                                                            .EMAC1_TXD3
		input  wire         hps_io_EMAC1_RX_CTL,                                                                     //                                                                            .EMAC1_RX_CTL
		output wire         hps_io_EMAC1_TX_CTL,                                                                     //                                                                            .EMAC1_TX_CTL
		input  wire         hps_io_EMAC1_RX_CLK,                                                                     //                                                                            .EMAC1_RX_CLK
		input  wire         hps_io_EMAC1_RXD0,                                                                       //                                                                            .EMAC1_RXD0
		input  wire         hps_io_EMAC1_RXD1,                                                                       //                                                                            .EMAC1_RXD1
		input  wire         hps_io_EMAC1_RXD2,                                                                       //                                                                            .EMAC1_RXD2
		input  wire         hps_io_EMAC1_RXD3,                                                                       //                                                                            .EMAC1_RXD3
		inout  wire         hps_io_EMAC1_MDIO,                                                                       //                                                                            .EMAC1_MDIO
		output wire         hps_io_EMAC1_MDC,                                                                        //                                                                            .EMAC1_MDC
		inout  wire         hps_io_SDMMC_CMD,                                                                        //                                                                            .SDMMC_CMD
		inout  wire         hps_io_SDMMC_D0,                                                                         //                                                                            .SDMMC_D0
		inout  wire         hps_io_SDMMC_D1,                                                                         //                                                                            .SDMMC_D1
		inout  wire         hps_io_SDMMC_D2,                                                                         //                                                                            .SDMMC_D2
		inout  wire         hps_io_SDMMC_D3,                                                                         //                                                                            .SDMMC_D3
		inout  wire         hps_io_SDMMC_D4,                                                                         //                                                                            .SDMMC_D4
		inout  wire         hps_io_SDMMC_D5,                                                                         //                                                                            .SDMMC_D5
		inout  wire         hps_io_SDMMC_D6,                                                                         //                                                                            .SDMMC_D6
		inout  wire         hps_io_SDMMC_D7,                                                                         //                                                                            .SDMMC_D7
		output wire         hps_io_SDMMC_CCLK,                                                                       //                                                                            .SDMMC_CCLK
		output wire         hps_io_SPIM0_CLK,                                                                        //                                                                            .SPIM0_CLK
		output wire         hps_io_SPIM0_MOSI,                                                                       //                                                                            .SPIM0_MOSI
		input  wire         hps_io_SPIM0_MISO,                                                                       //                                                                            .SPIM0_MISO
		output wire         hps_io_SPIM0_SS0_N,                                                                      //                                                                            .SPIM0_SS0_N
		output wire         hps_io_SPIM1_CLK,                                                                        //                                                                            .SPIM1_CLK
		output wire         hps_io_SPIM1_MOSI,                                                                       //                                                                            .SPIM1_MOSI
		input  wire         hps_io_SPIM1_MISO,                                                                       //                                                                            .SPIM1_MISO
		output wire         hps_io_SPIM1_SS0_N,                                                                      //                                                                            .SPIM1_SS0_N
		output wire         hps_io_SPIM1_SS1_N,                                                                      //                                                                            .SPIM1_SS1_N
		input  wire         hps_io_UART1_RX,                                                                         //                                                                            .UART1_RX
		output wire         hps_io_UART1_TX,                                                                         //                                                                            .UART1_TX
		inout  wire         hps_io_I2C1_SDA,                                                                         //                                                                            .I2C1_SDA
		inout  wire         hps_io_I2C1_SCL,                                                                         //                                                                            .I2C1_SCL
		input  wire         hps_io_hps_osc_clk,                                                                      //                                                                            .hps_osc_clk
		inout  wire         hps_io_gpio0_io11,                                                                       //                                                                            .gpio0_io11
		inout  wire         hps_io_gpio0_io12,                                                                       //                                                                            .gpio0_io12
		inout  wire         hps_io_gpio0_io13,                                                                       //                                                                            .gpio0_io13
		inout  wire         hps_io_gpio0_io14,                                                                       //                                                                            .gpio0_io14
		inout  wire         hps_io_gpio0_io15,                                                                       //                                                                            .gpio0_io15
		inout  wire         hps_io_gpio0_io16,                                                                       //                                                                            .gpio0_io16
		inout  wire         hps_io_gpio0_io17,                                                                       //                                                                            .gpio0_io17
		inout  wire         hps_io_gpio0_io18,                                                                       //                                                                            .gpio0_io18
		inout  wire         hps_io_gpio1_io16,                                                                       //                                                                            .gpio1_io16
		inout  wire         hps_io_gpio1_io17,                                                                       //                                                                            .gpio1_io17
		output wire         agilex_hps_h2f_reset_reset,                                                              //                                                        agilex_hps_h2f_reset.reset
		input  wire [31:0]  f2h_irq1_irq,                                                                            //                                                                    f2h_irq1.irq
		input  wire         emif_hps_pll_ref_clk_clk,                                                                //                                                        emif_hps_pll_ref_clk.clk
		input  wire         emif_hps_oct_oct_rzqin,                                                                  //                                                                emif_hps_oct.oct_rzqin
		output wire [0:0]   emif_hps_mem_mem_ck,                                                                     //                                                                emif_hps_mem.mem_ck
		output wire [0:0]   emif_hps_mem_mem_ck_n,                                                                   //                                                                            .mem_ck_n
		output wire [16:0]  emif_hps_mem_mem_a,                                                                      //                                                                            .mem_a
		output wire [0:0]   emif_hps_mem_mem_act_n,                                                                  //                                                                            .mem_act_n
		output wire [1:0]   emif_hps_mem_mem_ba,                                                                     //                                                                            .mem_ba
		output wire [0:0]   emif_hps_mem_mem_bg,                                                                     //                                                                            .mem_bg
		output wire [0:0]   emif_hps_mem_mem_cke,                                                                    //                                                                            .mem_cke
		output wire [1:0]   emif_hps_mem_mem_cs_n,                                                                   //                                                                            .mem_cs_n
		output wire [0:0]   emif_hps_mem_mem_odt,                                                                    //                                                                            .mem_odt
		output wire [0:0]   emif_hps_mem_mem_reset_n,                                                                //                                                                            .mem_reset_n
		output wire [0:0]   emif_hps_mem_mem_par,                                                                    //                                                                            .mem_par
		input  wire [0:0]   emif_hps_mem_mem_alert_n,                                                                //                                                                            .mem_alert_n
		inout  wire [8:0]   emif_hps_mem_mem_dqs,                                                                    //                                                                            .mem_dqs
		inout  wire [8:0]   emif_hps_mem_mem_dqs_n,                                                                  //                                                                            .mem_dqs_n
		inout  wire [71:0]  emif_hps_mem_mem_dq,                                                                     //                                                                            .mem_dq
		inout  wire [8:0]   emif_hps_mem_mem_dbi_n,                                                                  //                                                                            .mem_dbi_n
		output wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_rst_ack_n_export,                             //                        j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_rst_ack_n.export
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_txlclk_ctrl_export,                              //                         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_txlclk_ctrl.export
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_txfclk_ctrl_export,                              //                         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_txfclk_ctrl.export
		input  wire [511:0] j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avst_data,                                    //                             j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avst.data
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avst_valid,                                   //                                                                            .valid
		output wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avst_ready,                                   //                                                                            .ready
		input  wire [47:0]  j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_cmd_data,                                     //                              j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_cmd.data
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_cmd_valid,                                    //                                                                            .valid
		output wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_cmd_ready,                                    //                                                                            .ready
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_sysref_export,                                //                           j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_sysref.export
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rxlclk_ctrl_export,                              //                         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rxlclk_ctrl.export
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rxfclk_ctrl_export,                              //                         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rxfclk_ctrl.export
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_sysref_export,                                //                           j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_sysref.export
		output wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_rst_ack_n_export,                             //                        j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_rst_ack_n.export
		output wire [511:0] j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avst_data,                                    //                             j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avst.data
		output wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avst_valid,                                   //                                                                            .valid
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avst_ready,                                   //                                                                            .ready
		output wire [47:0]  j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_cmd_data,                                     //                              j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_cmd.data
		output wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_cmd_valid,                                    //                                                                            .valid
		input  wire         j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_cmd_ready,                                    //                                                                            .ready
		output wire [7:0]   j204c_f_rx_tx_ip_intel_jesd204c_f_tx_serial_data_export,                                 //                            j204c_f_rx_tx_ip_intel_jesd204c_f_tx_serial_data.export
		output wire [7:0]   j204c_f_rx_tx_ip_intel_jesd204c_f_tx_serial_data_n_export,                               //                          j204c_f_rx_tx_ip_intel_jesd204c_f_tx_serial_data_n.export
		input  wire [7:0]   j204c_f_rx_tx_ip_intel_jesd204c_f_rx_serial_data_export,                                 //                            j204c_f_rx_tx_ip_intel_jesd204c_f_rx_serial_data.export
		input  wire [7:0]   j204c_f_rx_tx_ip_intel_jesd204c_f_rx_serial_data_n_export,                               //                          j204c_f_rx_tx_ip_intel_jesd204c_f_rx_serial_data_n.export
		input  wire         j204c_f_rx_tx_ip_jesd_link_clk_in_clk_clk,                                               //                                       j204c_f_rx_tx_ip_jesd_link_clk_in_clk.clk
		output wire         j204c_f_rx_tx_ip_reset_out1_reset,                                                       //                                                 j204c_f_rx_tx_ip_reset_out1.reset
		output wire         j204c_f_rx_tx_ip_reset_out2_reset,                                                       //                                                 j204c_f_rx_tx_ip_reset_out2.reset
		output wire         j204c_f_rx_tx_ip_reset_out4_reset,                                                       //                                                 j204c_f_rx_tx_ip_reset_out4.reset
		input  wire         j204c_f_rx_tx_ip_reset1_dsrt_qual_reset1_dsrt_qual,                                      //                                           j204c_f_rx_tx_ip_reset1_dsrt_qual.reset1_dsrt_qual
		input  wire         j204c_f_rx_tx_ip_reset2_dsrt_qual_reset2_dsrt_qual,                                      //                                           j204c_f_rx_tx_ip_reset2_dsrt_qual.reset2_dsrt_qual
		input  wire         j204c_f_rx_tx_ip_reset4_dsrt_qual_reset4_dsrt_qual,                                      //                                           j204c_f_rx_tx_ip_reset4_dsrt_qual.reset4_dsrt_qual
		input  wire         j204c_f_rx_tx_ip_systemclk_f_refclk_fgt_in_refclk_fgt_0,                                 //                                     j204c_f_rx_tx_ip_systemclk_f_refclk_fgt.in_refclk_fgt_0
		input  wire [3:0]   button_pio_external_connection_export,                                                   //                                              button_pio_external_connection.export
		input  wire [3:0]   dipsw_pio_external_connection_export,                                                    //                                               dipsw_pio_external_connection.export
		input  wire [2:0]   led_pio_external_connection_in_port,                                                     //                                                 led_pio_external_connection.in_port
		output wire [2:0]   led_pio_external_connection_out_port,                                                    //                                                                            .out_port
		input  wire         ddc_avst_sink_avst_sink_valid,                                                           //                                                               ddc_avst_sink.avst_sink_valid
		input  wire [7:0]   ddc_avst_sink_avst_sink_channel,                                                         //                                                                            .avst_sink_channel
		input  wire [31:0]  ddc_avst_sink_avst_sink_data_l1,                                                         //                                                                            .avst_sink_data_l1
		input  wire [31:0]  ddc_avst_sink_avst_sink_data_l2,                                                         //                                                                            .avst_sink_data_l2
		input  wire [31:0]  ddc_avst_sink_avst_sink_data_l3,                                                         //                                                                            .avst_sink_data_l3
		input  wire [31:0]  ddc_avst_sink_avst_sink_data_l4,                                                         //                                                                            .avst_sink_data_l4
		input  wire [31:0]  ddc_avst_sink_avst_sink_data_l5,                                                         //                                                                            .avst_sink_data_l5
		input  wire [31:0]  ddc_avst_sink_avst_sink_data_l6,                                                         //                                                                            .avst_sink_data_l6
		input  wire [31:0]  ddc_avst_sink_avst_sink_data_l7,                                                         //                                                                            .avst_sink_data_l7
		input  wire [31:0]  ddc_avst_sink_avst_sink_data_l8,                                                         //                                                                            .avst_sink_data_l8
		output wire         duc_avst_source_duc_avst_source_valid,                                                   //                                                             duc_avst_source.duc_avst_source_valid
		output wire [31:0]  duc_avst_source_duc_avst_source_data0,                                                   //                                                                            .duc_avst_source_data0
		output wire [31:0]  duc_avst_source_duc_avst_source_data1,                                                   //                                                                            .duc_avst_source_data1
		output wire [31:0]  duc_avst_source_duc_avst_source_data2,                                                   //                                                                            .duc_avst_source_data2
		output wire [31:0]  duc_avst_source_duc_avst_source_data3,                                                   //                                                                            .duc_avst_source_data3
		output wire [31:0]  duc_avst_source_duc_avst_source_data4,                                                   //                                                                            .duc_avst_source_data4
		output wire [31:0]  duc_avst_source_duc_avst_source_data5,                                                   //                                                                            .duc_avst_source_data5
		output wire [31:0]  duc_avst_source_duc_avst_source_data6,                                                   //                                                                            .duc_avst_source_data6
		output wire [31:0]  duc_avst_source_duc_avst_source_data7,                                                   //                                                                            .duc_avst_source_data7
		output wire [7:0]   duc_avst_source_duc_avst_source_channel,                                                 //                                                                            .duc_avst_source_channel
		input  wire         avst_tx_ptp_i_av_st_tx_skip_crc,                                                         //                                                                 avst_tx_ptp.i_av_st_tx_skip_crc
		input  wire [1:0]   avst_tx_ptp_i_av_st_tx_ptp_ts_valid,                                                     //                                                                            .i_av_st_tx_ptp_ts_valid
		input  wire         avst_tx_ptp_i_av_st_tx_ptp_ins_ets,                                                      //                                                                            .i_av_st_tx_ptp_ins_ets
		input  wire         avst_tx_ptp_i_av_st_tx_ptp_ins_cf,                                                       //                                                                            .i_av_st_tx_ptp_ins_cf
		input  wire [95:0]  avst_tx_ptp_i_av_st_tx_ptp_tx_its,                                                       //                                                                            .i_av_st_tx_ptp_tx_its
		input  wire [6:0]   avst_tx_ptp_i_av_st_tx_ptp_asym_p2p_idx,                                                 //                                                                            .i_av_st_tx_ptp_asym_p2p_idx
		input  wire         avst_tx_ptp_i_av_st_tx_ptp_asym_sign,                                                    //                                                                            .i_av_st_tx_ptp_asym_sign
		input  wire         avst_tx_ptp_i_av_st_tx_ptp_asym,                                                         //                                                                            .i_av_st_tx_ptp_asym
		input  wire         avst_tx_ptp_i_av_st_tx_ptp_p2p,                                                          //                                                                            .i_av_st_tx_ptp_p2p
		input  wire         avst_tx_ptp_i_av_st_tx_ptp_ts_format,                                                    //                                                                            .i_av_st_tx_ptp_ts_format
		input  wire         avst_tx_ptp_i_av_st_tx_ptp_update_eb,                                                    //                                                                            .i_av_st_tx_ptp_update_eb
		input  wire         avst_tx_ptp_i_av_st_tx_ptp_zero_csum,                                                    //                                                                            .i_av_st_tx_ptp_zero_csum
		input  wire [15:0]  avst_tx_ptp_i_av_st_tx_ptp_eb_offset,                                                    //                                                                            .i_av_st_tx_ptp_eb_offset
		input  wire [15:0]  avst_tx_ptp_i_av_st_tx_ptp_csum_offset,                                                  //                                                                            .i_av_st_tx_ptp_csum_offset
		input  wire [15:0]  avst_tx_ptp_i_av_st_tx_ptp_cf_offset,                                                    //                                                                            .i_av_st_tx_ptp_cf_offset
		input  wire [15:0]  avst_tx_ptp_i_av_st_tx_ptp_ts_offset,                                                    //                                                                            .i_av_st_tx_ptp_ts_offset
		input  wire         avst_axist_bridge_0_axit_tx_if_tready,                                                   //                                              avst_axist_bridge_0_axit_tx_if.tready
		output wire         avst_axist_bridge_0_axit_tx_if_tvalid,                                                   //                                                                            .tvalid
		output wire [63:0]  avst_axist_bridge_0_axit_tx_if_tdata,                                                    //                                                                            .tdata
		output wire         avst_axist_bridge_0_axit_tx_if_tlast,                                                    //                                                                            .tlast
		output wire [7:0]   avst_axist_bridge_0_axit_tx_if_tkeep,                                                    //                                                                            .tkeep
		output wire [1:0]   avst_axist_bridge_0_axit_tx_if_tuser,                                                    //                                                                            .tuser
		output wire [93:0]  axist_tx_user_o_axi_st_tx_tuser_ptp,                                                     //                                                               axist_tx_user.o_axi_st_tx_tuser_ptp
		output wire [327:0] axist_tx_user_o_axi_st_tx_tuser_ptp_extended,                                            //                                                                            .o_axi_st_tx_tuser_ptp_extended
		output wire [39:0]  avst_rx_ptp_o_av_st_rxstatus_data,                                                       //                                                                 avst_rx_ptp.o_av_st_rxstatus_data
		output wire         avst_rx_ptp_o_av_st_rxstatus_valid,                                                      //                                                                            .o_av_st_rxstatus_valid
		output wire [95:0]  avst_rx_ptp_o_av_st_ptp_rx_its,                                                          //                                                                            .o_av_st_ptp_rx_its
		input  wire [4:0]   axist_rx_user_i_axi_st_rx_tuser_sts,                                                     //                                                               axist_rx_user.i_axi_st_rx_tuser_sts
		input  wire [31:0]  axist_rx_user_i_axi_st_rx_tuser_sts_extended,                                            //                                                                            .i_axi_st_rx_tuser_sts_extended
		input  wire [95:0]  axist_rx_user_i_axi_st_rx_ingrts0_tdata,                                                 //                                                                            .i_axi_st_rx_ingrts0_tdata
		input  wire         axist_rx_user_i_axi_st_rx_ingrts0_tvalid,                                                //                                                                            .i_axi_st_rx_ingrts0_tvalid
		output wire [21:0]  ptp_tod_concat_out_o_mac_ptp_fp,                                                         //                                                          ptp_tod_concat_out.o_mac_ptp_fp
		output wire         ptp_tod_concat_out_o_mac_ptp_ts_req,                                                     //                                                                            .o_mac_ptp_ts_req
		input  wire         ptp_tod_concat_out_i_mac_ptp_tx_ets_valid,                                               //                                                                            .i_mac_ptp_tx_ets_valid
		input  wire [95:0]  ptp_tod_concat_out_i_mac_ptp_tx_ets,                                                     //                                                                            .i_mac_ptp_tx_ets
		input  wire [21:0]  ptp_tod_concat_out_i_mac_ptp_tx_ets_fp,                                                  //                                                                            .i_mac_ptp_tx_ets_fp
		input  wire         ptp_tod_concat_out_i_mac_ptp_rx_its_valid,                                               //                                                                            .i_mac_ptp_rx_its_valid
		input  wire [95:0]  ptp_tod_concat_out_i_mac_ptp_rx_its,                                                     //                                                                            .i_mac_ptp_rx_its
		input  wire [19:0]  ptp_tod_concat_out_i_ext_ptp_fp,                                                         //                                                                            .i_ext_ptp_fp
		input  wire         ptp_tod_concat_out_i_ext_ptp_ts_req,                                                     //                                                                            .i_ext_ptp_ts_req
		output wire         ptp_tod_concat_out_o_ext_ptp_tx_ets_valid,                                               //                                                                            .o_ext_ptp_tx_ets_valid
		output wire [95:0]  ptp_tod_concat_out_o_ext_ptp_tx_ets,                                                     //                                                                            .o_ext_ptp_tx_ets
		output wire [19:0]  ptp_tod_concat_out_o_ext_ptp_tx_ets_fp,                                                  //                                                                            .o_ext_ptp_tx_ets_fp
		output wire [95:0]  ptp_tod_concat_out_o_ext_ptp_rx_its,                                                     //                                                                            .o_ext_ptp_rx_its
		output wire         ptp_tod_concat_out_o_ext_ptp_rx_its_valid,                                               //                                                                            .o_ext_ptp_rx_its_valid
		input  wire         phipps_peak_0_rx_pcs_ready_rx_pcs_ready,                                                 //                                                  phipps_peak_0_rx_pcs_ready.rx_pcs_ready
		input  wire         phipps_peak_0_tx_lanes_stable_tx_lanes_stable,                                           //                                               phipps_peak_0_tx_lanes_stable.tx_lanes_stable
		output wire         phipps_peak_0_lphy_ss_top_0_lphy_ss_top_duc_ddc_lpbk_en_data,                            //                     phipps_peak_0_lphy_ss_top_0_lphy_ss_top_duc_ddc_lpbk_en.data
		input  wire         rst_dsp_in_reset_reset,                                                                  //                                                            rst_dsp_in_reset.reset
		input  wire         rst_eth_in_reset_reset,                                                                  //                                                            rst_eth_in_reset.reset
		input  wire         rst_csr_act_high_in_reset_reset,                                                         //                                                   rst_csr_act_high_in_reset.reset
		input  wire         rst_csr_in_reset_reset_n,                                                                //                                                            rst_csr_in_reset.reset_n
		input  wire         clk_100_clk,                                                                             //                                                                     clk_100.clk
		input  wire         dma_subsys_port0_rx_dma_resetn_reset_n,                                                  //                                      dma_subsys_port0_rx_dma_resetn_reset_n.reset_n
		input  wire         dma_subsys_port1_rx_dma_resetn_reset_n,                                                  //                                      dma_subsys_port1_rx_dma_resetn_reset_n.reset_n
		input  wire         qsys_top_master_todclk_0_in_clk_clk,                                                     //                                             qsys_top_master_todclk_0_in_clk.clk
		input  wire         reset_reset_n,                                                                           //                                                                       reset.reset_n
		output wire         ninit_done_ninit_done,                                                                   //                                                                  ninit_done.ninit_done
		input  wire         tod_timestamp_96b_0_pps_in_pps_in,                                                       //                                                  tod_timestamp_96b_0_pps_in.pps_in
		output wire         master_tod_top_0_pulse_per_second_pps,                                                   //                                           master_tod_top_0_pulse_per_second.pps
		input  wire         mtod_subsys_master_tod_top_0_i_upstr_pll_lock,                                           //                                    mtod_subsys_master_tod_top_0_i_upstr_pll.lock
		input  wire         mtod_subsys_pps_in_pulse_per_second,                                                     //                                                          mtod_subsys_pps_in.pulse_per_second
		input  wire         tod_slave_subsys_oran_tod_stack_tx_pll_locked_lock,                                      //                               tod_slave_subsys_oran_tod_stack_tx_pll_locked.lock
		input  wire         tod_slave_subsys_port_8_tod_stack_tx_pll_locked_lock                                     //                             tod_slave_subsys_port_8_tod_stack_tx_pll_locked.lock
	);

	wire          dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid;          // dma_subsys:dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid -> phipps_peak_0:ecpri_ext_sink_valid
	wire   [63:0] dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data;           // dma_subsys:dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data -> phipps_peak_0:ecpri_ext_sink_data
	wire          dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready;          // phipps_peak_0:ecpri_ext_sink_ready -> dma_subsys:dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready
	wire          dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket;  // dma_subsys:dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket -> phipps_peak_0:ecpri_ext_sink_startofpacket
	wire          dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket;    // dma_subsys:dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket -> phipps_peak_0:ecpri_ext_sink_endofpacket
	wire    [0:0] dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error;          // dma_subsys:dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error -> phipps_peak_0:ecpri_ext_sink_error
	wire    [2:0] dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty;          // dma_subsys:dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty -> phipps_peak_0:ecpri_ext_sink_empty
	wire          phipps_peak_0_dxc_avst_selctd_cap_intf_valid;                                           // phipps_peak_0:dxc_avst_selctd_cap_intf_valid -> dfd_subsystem:dxc_avst_sink_dsp_capture_valid
	wire   [31:0] phipps_peak_0_dxc_avst_selctd_cap_intf_data;                                            // phipps_peak_0:dxc_avst_selctd_cap_intf_data -> dfd_subsystem:dxc_avst_sink_dsp_capture_data
	wire    [2:0] phipps_peak_0_dxc_avst_selctd_cap_intf_channel;                                         // phipps_peak_0:dxc_avst_selctd_cap_intf_channel -> dfd_subsystem:dxc_avst_sink_dsp_capture_channel
	wire          phipps_peak_0_ecpri_ext_source_valid;                                                   // phipps_peak_0:ecpri_ext_source_valid -> dma_subsys:dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_valid
	wire   [63:0] phipps_peak_0_ecpri_ext_source_data;                                                    // phipps_peak_0:ecpri_ext_source_data -> dma_subsys:dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_data
	wire          phipps_peak_0_ecpri_ext_source_startofpacket;                                           // phipps_peak_0:ecpri_ext_source_startofpacket -> dma_subsys:dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_startofpacket
	wire          phipps_peak_0_ecpri_ext_source_endofpacket;                                             // phipps_peak_0:ecpri_ext_source_endofpacket -> dma_subsys:dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_endofpacket
	wire    [5:0] phipps_peak_0_ecpri_ext_source_error;                                                   // phipps_peak_0:ecpri_ext_source_error -> dma_subsys:dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_error
	wire    [2:0] phipps_peak_0_ecpri_ext_source_empty;                                                   // phipps_peak_0:ecpri_ext_source_empty -> dma_subsys:dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_empty
	wire          phipps_peak_0_lphy_avst_selctd_cap_intf_valid;                                          // phipps_peak_0:lphy_avst_selctd_cap_intf_valid -> dfd_subsystem:lphy_avst_sink_dsp_capture_valid
	wire   [31:0] phipps_peak_0_lphy_avst_selctd_cap_intf_data;                                           // phipps_peak_0:lphy_avst_selctd_cap_intf_data -> dfd_subsystem:lphy_avst_sink_dsp_capture_data
	wire    [2:0] phipps_peak_0_lphy_avst_selctd_cap_intf_channel;                                        // phipps_peak_0:lphy_avst_selctd_cap_intf_channel -> dfd_subsystem:lphy_avst_sink_dsp_capture_channel
	wire          hssi_ss_1_p0_axi_st_rx_interface_tvalid;                                                // hssi_ss_1:p0_ss_app_st_rx_tvalid -> phipps_peak_0:avst_axist_bridge_0_axist_rx_if_tvalid
	wire    [6:0] hssi_ss_1_p0_axi_st_rx_interface_tuser;                                                 // hssi_ss_1:p0_ss_app_st_rx_tuser_client -> phipps_peak_0:avst_axist_bridge_0_axist_rx_if_tuser
	wire    [7:0] hssi_ss_1_p0_axi_st_rx_interface_tkeep;                                                 // hssi_ss_1:p0_ss_app_st_rx_tkeep -> phipps_peak_0:avst_axist_bridge_0_axist_rx_if_tkeep
	wire   [63:0] hssi_ss_1_p0_axi_st_rx_interface_tdata;                                                 // hssi_ss_1:p0_ss_app_st_rx_tdata -> phipps_peak_0:avst_axist_bridge_0_axist_rx_if_tdata
	wire          hssi_ss_1_p0_axi_st_rx_interface_tlast;                                                 // hssi_ss_1:p0_ss_app_st_rx_tlast -> phipps_peak_0:avst_axist_bridge_0_axist_rx_if_tlast
	wire          dma_subsys_acp_bridge_in_clk_clk;                                                       // dma_subsys:acp_bridge_in_clk_clk -> [hps_sub_sys:acp_0_clock_clk, mm_interconnect_2:dma_subsys_acp_bridge_in_clk_clk, rst_controller_001:clk, rst_controller_008:clk]
	wire          sys_manager_clk_100_out_clk_clk;                                                        // sys_manager:clk_100_out_clk_clk -> [dma_subsys:dma_clk_100_in_clk_clk, ftile_debug_status_pio_0:clk, hps_sub_sys:acp_0_csr_clock_clk, hps_sub_sys:agilex_hps_h2f_axi_clock_clk, hps_sub_sys:agilex_hps_h2f_lw_axi_clock_clk, hssi_ss_1:app_ss_lite_clk, irq_mapper_001:clk, j204c_f_rx_tx_ip:mgmt_clk_in_clk_clk, jtg_mst:clk_clk, mm_interconnect_0:sys_manager_clk_100_out_clk_clk, mm_interconnect_1:sys_manager_clk_100_out_clk_clk, mm_interconnect_2:sys_manager_clk_100_out_clk_clk, mm_interconnect_3:sys_manager_clk_100_out_clk_clk, ocm:clk, periph:clk_clk, qsfpdd_status_pio:clk, rst_controller:clk, rst_controller_002:clk, sys_ctrl_pio_0:clk, sys_manager:dma_subsys_port0_rx_dma_resetn_clk_clk, sys_manager:dma_subsys_port1_rx_dma_resetn_clk_clk, sys_manager:ftile_iopll_ptp_sampling_refclk_clk, sys_manager:rst_in_clk_clk, sys_manager:sysid_clk_clk, tod_subsys_0:mtod_subsys_clk100_in_clk_clk, tod_subsys_0:tod_slave_tod_subsys_clk_100_in_clk_clk]
	wire          clk_ss_0_clk_csr_out_clk_clk;                                                           // clk_ss_0:clk_csr_out_clk_clk -> [dfd_subsystem:clock_csr_clk, mm_interconnect_0:clk_ss_0_clk_csr_out_clk_clk, mm_interconnect_1:clk_ss_0_clk_csr_out_clk_clk, phipps_peak_0:clock_bridge_csr_in_clk_clk, rst_controller_006:clk, rst_ss_0:reset_bridge_act_high_clk_clk, rst_ss_0:rst_csr_clk_clk, tod_subsys_0:clock_bridge_100_in_clk_clk]
	wire          clk_ss_0_clk_dsp_out_clk_clk;                                                           // clk_ss_0:clk_dsp_out_clk_clk -> [dfd_subsystem:dsp_in_clk_clk, phipps_peak_0:clock_bridge_dsp_in_clk_clk, rst_ss_0:dsp_rst_cntrl_clk_clk]
	wire          clk_ss_0_clk_eth_out_clk_clk;                                                           // clk_ss_0:clk_eth_out_clk_clk -> [dfd_subsystem:eth_in_clk_clk, phipps_peak_0:clock_bridge_eth_in_clk_clk, rst_ss_0:eth_rst_cntrl_clk_clk]
	wire          clk_ss_0_clk_ftile_402_out_clk_clk;                                                     // clk_ss_0:clk_ftile_402_out_clk_clk -> [dma_subsys:dma_subsys_port8_ts_chs_compl_0_clk_bus_in_clk, dma_subsys:oclk_pll_port8_in_clk_clk, hssi_ss_1:p0_app_ss_st_rx_clk, hssi_ss_1:p0_app_ss_st_tx_clk, phipps_peak_0:clock_bridge_ecpri_rx_in_clk_clk, phipps_peak_0:clock_bridge_ecpri_tx_in_clk_clk, rst_ss_0:ecpri_rst_cntrl_clk_clk, tod_subsys_0:cdc_pipeline_0_dst_clk_clk]
	wire          dma_subsys_dma_clk_out_bridge_0_out_clk_clk;                                            // dma_subsys:dma_clk_out_bridge_0_out_clk_clk -> [hps_sub_sys:agilex_hps_f2h_axi_clock_clk, mm_interconnect_2:dma_subsys_dma_clk_out_bridge_0_out_clk_clk, rst_controller_007:clk]
	wire          sys_manager_ftile_iopll_ptp_sampling_outclk0_clk;                                       // sys_manager:ftile_iopll_ptp_sampling_outclk0_clk -> hssi_ss_1:i_p0_clk_ptp_sample
	wire          sys_manager_ftile_iopll_todsync_sampling_outclk0_clk;                                   // sys_manager:ftile_iopll_todsync_sampling_outclk0_clk -> [tod_subsys_0:tod_slave_oran_tod_stack_todsync_sample_clk_clk, tod_subsys_0:tod_slave_port_8_tod_stack_todsync_sample_clk_clk]
	wire          hssi_ss_1_o_p0_clk_pll_clk;                                                             // hssi_ss_1:o_p0_clk_pll -> [clk_ss_0:clk_ftile_402_in_clk_clk, clk_ss_0:ftile_in_clk_clk]
	wire          hssi_ss_1_o_p0_clk_rec_div_clk_signal;                                                  // hssi_ss_1:o_p0_clk_rec_div -> [clk_ss_0:clk_eth_in_clk_clk, clk_ss_0:clock_bridge_rec_rx_in_clk_clk, hssi_ss_1:i_p0_clk_rx_tod, rst_controller_003:clk, rst_ss_0:reset_bridge_rec_rx_clk_clk, tod_subsys_0:tod_slave_oran_tod_stack_rx_clk_clk, tod_subsys_0:tod_slave_port_8_tod_stack_rx_clk_clk]
	wire          hssi_ss_1_o_p0_clk_tx_div_clk;                                                          // hssi_ss_1:o_p0_clk_tx_div -> [hssi_ss_1:i_p0_clk_tx_tod, rst_controller_004:clk, rst_ss_0:reset_bridge_tx_div_clk_clk, tod_subsys_0:tod_slave_oran_tod_stack_tx_clk_clk, tod_subsys_0:tod_slave_port_8_tod_stack_tx_clk_clk]
	wire          sys_manager_qsys_top_master_todclk_0_out_clk_clk;                                       // sys_manager:qsys_top_master_todclk_0_out_clk_clk -> [rst_controller_005:clk, sys_manager:ftile_iopll_todsync_sampling_refclk_clk, tod_subsys_0:clock_bridge_156_in_clk_clk, tod_subsys_0:mtod_subsys_pps_load_tod_0_period_clock_clk, tod_subsys_0:tod_slave_tod_subsys_mtod_clk_in_clk_clk]
	wire   [55:0] phipps_peak_0_radio_config_status_dup2_radio_config_status;                             // phipps_peak_0:radio_config_status_dup2_radio_config_status -> dfd_subsystem:capture_if_radio_config_status_radio_config_status
	wire          phipps_peak_0_rst_soft_n_dup4_rst_soft_n;                                               // phipps_peak_0:rst_soft_n_dup4_rst_soft_n -> dfd_subsystem:capture_if_reset_soft_n_rst_soft_n
	wire   [95:0] tod_subsys_0_cdc_pipeline_0_dataout_data;                                               // tod_subsys_0:cdc_pipeline_0_dataout_data -> phipps_peak_0:xran_timestamp_tod_in_data
	wire          tod_subsys_0_tod_timestamp_96b_0_rfp_sync_pul_data;                                     // tod_subsys_0:tod_timestamp_96b_0_rfp_sync_pul_data -> phipps_peak_0:dxc_ss_top_0_rfp_pulse_data
	wire          sys_manager_ftile_iopll_todsync_sampling_locked_lock;                                   // sys_manager:ftile_iopll_todsync_sampling_locked_lock -> tod_subsys_0:tod_slave_todsync_sample_plllock_split_conduit_end_lock
	wire   [31:0] dfd_subsystem_interface_sel_data;                                                       // dfd_subsystem:interface_sel_data -> phipps_peak_0:interface_sel_data
	wire          tod_subsys_0_tod_timestamp_96b_0_rfp_sync_pul_dup_data;                                 // tod_subsys_0:tod_timestamp_96b_0_rfp_sync_pul_dup_data -> phipps_peak_0:lphy_ss_top_0_frame_status_counter_reset_data
	wire          tod_subsys_0_tod_slave_port_8_tod_stack_rx_tod_interface_tvalid;                        // tod_subsys_0:tod_slave_port_8_tod_stack_rx_tod_interface_tvalid -> hssi_ss_1:p0_app_ss_st_rxtod_tvalid
	wire   [95:0] tod_subsys_0_tod_slave_port_8_tod_stack_rx_tod_interface_tdata;                         // tod_subsys_0:tod_slave_port_8_tod_stack_rx_tod_interface_tdata -> hssi_ss_1:p0_app_ss_st_rxtod_tdata
	wire          tod_subsys_0_tod_slave_port_8_tod_stack_tx_tod_interface_tvalid;                        // tod_subsys_0:tod_slave_port_8_tod_stack_tx_tod_interface_tvalid -> hssi_ss_1:p0_app_ss_st_txtod_tvalid
	wire   [95:0] tod_subsys_0_tod_slave_port_8_tod_stack_tx_tod_interface_tdata;                         // tod_subsys_0:tod_slave_port_8_tod_stack_tx_tod_interface_tdata -> hssi_ss_1:p0_app_ss_st_txtod_tdata
	wire          tod_subsys_0_rx_oran_tod_time_of_day_96b_tvalid;                                        // tod_subsys_0:rx_oran_tod_time_of_day_96b_tvalid -> phipps_peak_0:ecpri_oran_top_0_oran_rx_tod_96b_data_tvalid
	wire   [95:0] tod_subsys_0_rx_oran_tod_time_of_day_96b_tdata;                                         // tod_subsys_0:rx_oran_tod_time_of_day_96b_tdata -> phipps_peak_0:ecpri_oran_top_0_oran_rx_tod_96b_data_tdata
	wire          tod_subsys_0_tx_oran_tod_time_of_day_96b_tvalid;                                        // tod_subsys_0:tx_oran_tod_time_of_day_96b_tvalid -> phipps_peak_0:ecpri_oran_top_0_oran_tx_tod_96b_data_tvalid
	wire   [95:0] tod_subsys_0_tx_oran_tod_time_of_day_96b_tdata;                                         // tod_subsys_0:tx_oran_tod_time_of_day_96b_tdata -> phipps_peak_0:ecpri_oran_top_0_oran_tx_tod_96b_data_tdata
	wire          sys_manager_dma_subsys_port0_rx_dma_resetn_out_reset_reset;                             // sys_manager:dma_subsys_port0_rx_dma_resetn_out_reset_reset_n -> dma_subsys:rx_dma_reset_bridge_0_in_reset_reset_n
	wire          sys_manager_dma_subsys_port1_rx_dma_resetn_out_reset_reset;                             // sys_manager:dma_subsys_port1_rx_dma_resetn_out_reset_reset_n -> dma_subsys:rx_dma_reset_bridge_1_in_reset_reset_n
	wire          rst_ss_0_dsp_rst_cntrl_reset_out_reset;                                                 // rst_ss_0:dsp_rst_cntrl_reset_out_reset -> [dfd_subsystem:dsp_in_reset_reset_n, phipps_peak_0:dsp_in_reset_reset_n]
	wire          rst_ss_0_ecpri_rst_cntrl_reset_out_reset;                                               // rst_ss_0:ecpri_rst_cntrl_reset_out_reset -> phipps_peak_0:rst_ecpri_n_reset_n
	wire          rst_ss_0_eth_rst_cntrl_reset_out_reset;                                                 // rst_ss_0:eth_rst_cntrl_reset_out_reset -> [dfd_subsystem:eth_in_reset_reset_n, phipps_peak_0:eth_in_reset_reset_n, tod_subsys_0:cdc_pipeline_0_rst_dst_clk_n_reset_n]
	wire          hssi_ss_1_o_p0_ereset_n_reset;                                                          // hssi_ss_1:o_p0_ereset_n -> rst_ss_0:ecpri_rst_cntrl_reset_in0_reset
	wire          rst_ss_0_rst_csr_out_reset_reset;                                                       // rst_ss_0:rst_csr_out_reset_reset_n -> [dfd_subsystem:reset_csr_reset_n, phipps_peak_0:csr_in_reset_reset_n, rst_controller_006:reset_in0, tod_subsys_0:reset_bridge_100_in_reset_reset_n]
	wire          sys_manager_rst_in_out_reset_reset;                                                     // sys_manager:rst_in_out_reset_reset_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_007:reset_in0, rst_controller_008:reset_in0, sys_manager:ftile_iopll_ptp_sampling_reset_reset, sys_manager:ftile_iopll_todsync_sampling_reset_reset]
	wire          dma_subsys_subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset_reset;                     // dma_subsys:subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset_reset_n -> hps_sub_sys:agilex_hps_f2h_axi_reset_reset_n
	wire    [1:0] hps_sub_sys_agilex_hps_h2f_axi_master_awburst;                                          // hps_sub_sys:agilex_hps_h2f_axi_master_awburst -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awburst
	wire    [7:0] hps_sub_sys_agilex_hps_h2f_axi_master_arlen;                                            // hps_sub_sys:agilex_hps_h2f_axi_master_arlen -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arlen
	wire   [15:0] hps_sub_sys_agilex_hps_h2f_axi_master_wstrb;                                            // hps_sub_sys:agilex_hps_h2f_axi_master_wstrb -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_wstrb
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_wready;                                           // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_wready -> hps_sub_sys:agilex_hps_h2f_axi_master_wready
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_axi_master_rid;                                              // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_rid -> hps_sub_sys:agilex_hps_h2f_axi_master_rid
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_rready;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_rready -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_rready
	wire    [7:0] hps_sub_sys_agilex_hps_h2f_axi_master_awlen;                                            // hps_sub_sys:agilex_hps_h2f_axi_master_awlen -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awlen
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_axi_master_arcache;                                          // hps_sub_sys:agilex_hps_h2f_axi_master_arcache -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arcache
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_wvalid;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_wvalid -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_wvalid
	wire   [31:0] hps_sub_sys_agilex_hps_h2f_axi_master_araddr;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_araddr -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_araddr
	wire    [2:0] hps_sub_sys_agilex_hps_h2f_axi_master_arprot;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_arprot -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arprot
	wire    [2:0] hps_sub_sys_agilex_hps_h2f_axi_master_awprot;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_awprot -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awprot
	wire  [127:0] hps_sub_sys_agilex_hps_h2f_axi_master_wdata;                                            // hps_sub_sys:agilex_hps_h2f_axi_master_wdata -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_wdata
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_arvalid;                                          // hps_sub_sys:agilex_hps_h2f_axi_master_arvalid -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arvalid
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_axi_master_awcache;                                          // hps_sub_sys:agilex_hps_h2f_axi_master_awcache -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awcache
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_axi_master_arid;                                             // hps_sub_sys:agilex_hps_h2f_axi_master_arid -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arid
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_arlock;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_arlock -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arlock
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_awlock;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_awlock -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awlock
	wire   [31:0] hps_sub_sys_agilex_hps_h2f_axi_master_awaddr;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_awaddr -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awaddr
	wire    [1:0] hps_sub_sys_agilex_hps_h2f_axi_master_bresp;                                            // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_bresp -> hps_sub_sys:agilex_hps_h2f_axi_master_bresp
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_arready;                                          // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arready -> hps_sub_sys:agilex_hps_h2f_axi_master_arready
	wire  [127:0] hps_sub_sys_agilex_hps_h2f_axi_master_rdata;                                            // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_rdata -> hps_sub_sys:agilex_hps_h2f_axi_master_rdata
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_awready;                                          // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awready -> hps_sub_sys:agilex_hps_h2f_axi_master_awready
	wire    [1:0] hps_sub_sys_agilex_hps_h2f_axi_master_arburst;                                          // hps_sub_sys:agilex_hps_h2f_axi_master_arburst -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arburst
	wire    [2:0] hps_sub_sys_agilex_hps_h2f_axi_master_arsize;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_arsize -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_arsize
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_bready;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_bready -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_bready
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_rlast;                                            // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_rlast -> hps_sub_sys:agilex_hps_h2f_axi_master_rlast
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_wlast;                                            // hps_sub_sys:agilex_hps_h2f_axi_master_wlast -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_wlast
	wire    [1:0] hps_sub_sys_agilex_hps_h2f_axi_master_rresp;                                            // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_rresp -> hps_sub_sys:agilex_hps_h2f_axi_master_rresp
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_axi_master_awid;                                             // hps_sub_sys:agilex_hps_h2f_axi_master_awid -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awid
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_axi_master_bid;                                              // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_bid -> hps_sub_sys:agilex_hps_h2f_axi_master_bid
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_bvalid;                                           // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_bvalid -> hps_sub_sys:agilex_hps_h2f_axi_master_bvalid
	wire    [2:0] hps_sub_sys_agilex_hps_h2f_axi_master_awsize;                                           // hps_sub_sys:agilex_hps_h2f_axi_master_awsize -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awsize
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_awvalid;                                          // hps_sub_sys:agilex_hps_h2f_axi_master_awvalid -> mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_awvalid
	wire          hps_sub_sys_agilex_hps_h2f_axi_master_rvalid;                                           // mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_master_rvalid -> hps_sub_sys:agilex_hps_h2f_axi_master_rvalid
	wire          jtg_mst_fpga_m2ocm_pb_m0_waitrequest;                                                   // mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_waitrequest -> jtg_mst:fpga_m2ocm_pb_m0_waitrequest
	wire  [127:0] jtg_mst_fpga_m2ocm_pb_m0_readdata;                                                      // mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_readdata -> jtg_mst:fpga_m2ocm_pb_m0_readdata
	wire          jtg_mst_fpga_m2ocm_pb_m0_debugaccess;                                                   // jtg_mst:fpga_m2ocm_pb_m0_debugaccess -> mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_debugaccess
	wire   [17:0] jtg_mst_fpga_m2ocm_pb_m0_address;                                                       // jtg_mst:fpga_m2ocm_pb_m0_address -> mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_address
	wire          jtg_mst_fpga_m2ocm_pb_m0_read;                                                          // jtg_mst:fpga_m2ocm_pb_m0_read -> mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_read
	wire   [15:0] jtg_mst_fpga_m2ocm_pb_m0_byteenable;                                                    // jtg_mst:fpga_m2ocm_pb_m0_byteenable -> mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_byteenable
	wire          jtg_mst_fpga_m2ocm_pb_m0_readdatavalid;                                                 // mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_readdatavalid -> jtg_mst:fpga_m2ocm_pb_m0_readdatavalid
	wire  [127:0] jtg_mst_fpga_m2ocm_pb_m0_writedata;                                                     // jtg_mst:fpga_m2ocm_pb_m0_writedata -> mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_writedata
	wire          jtg_mst_fpga_m2ocm_pb_m0_write;                                                         // jtg_mst:fpga_m2ocm_pb_m0_write -> mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_write
	wire    [0:0] jtg_mst_fpga_m2ocm_pb_m0_burstcount;                                                    // jtg_mst:fpga_m2ocm_pb_m0_burstcount -> mm_interconnect_0:jtg_mst_fpga_m2ocm_pb_m0_burstcount
	wire   [25:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awaddr;                                 // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_awaddr -> hssi_ss_1:app_ss_lite_awaddr
	wire    [1:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bresp;                                  // hssi_ss_1:ss_app_lite_bresp -> mm_interconnect_0:hssi_ss_1_axi4_lite_interface_bresp
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arready;                                // hssi_ss_1:ss_app_lite_arready -> mm_interconnect_0:hssi_ss_1_axi4_lite_interface_arready
	wire   [31:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rdata;                                  // hssi_ss_1:ss_app_lite_rdata -> mm_interconnect_0:hssi_ss_1_axi4_lite_interface_rdata
	wire    [3:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wstrb;                                  // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_wstrb -> hssi_ss_1:app_ss_lite_wstrb
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wready;                                 // hssi_ss_1:ss_app_lite_wready -> mm_interconnect_0:hssi_ss_1_axi4_lite_interface_wready
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awready;                                // hssi_ss_1:ss_app_lite_awready -> mm_interconnect_0:hssi_ss_1_axi4_lite_interface_awready
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rready;                                 // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_rready -> hssi_ss_1:app_ss_lite_rready
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bready;                                 // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_bready -> hssi_ss_1:app_ss_lite_bready
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wvalid;                                 // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_wvalid -> hssi_ss_1:app_ss_lite_wvalid
	wire   [25:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_araddr;                                 // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_araddr -> hssi_ss_1:app_ss_lite_araddr
	wire    [2:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arprot;                                 // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_arprot -> hssi_ss_1:app_ss_lite_arprot
	wire    [1:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rresp;                                  // hssi_ss_1:ss_app_lite_rresp -> mm_interconnect_0:hssi_ss_1_axi4_lite_interface_rresp
	wire    [2:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awprot;                                 // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_awprot -> hssi_ss_1:app_ss_lite_awprot
	wire   [31:0] mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wdata;                                  // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_wdata -> hssi_ss_1:app_ss_lite_wdata
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arvalid;                                // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_arvalid -> hssi_ss_1:app_ss_lite_arvalid
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bvalid;                                 // hssi_ss_1:ss_app_lite_bvalid -> mm_interconnect_0:hssi_ss_1_axi4_lite_interface_bvalid
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awvalid;                                // mm_interconnect_0:hssi_ss_1_axi4_lite_interface_awvalid -> hssi_ss_1:app_ss_lite_awvalid
	wire          mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rvalid;                                 // hssi_ss_1:ss_app_lite_rvalid -> mm_interconnect_0:hssi_ss_1_axi4_lite_interface_rvalid
	wire   [31:0] mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_readdata;                             // dma_subsys:dma_subsys_port8_csr_readdata -> mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_readdata
	wire          mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_waitrequest;                          // dma_subsys:dma_subsys_port8_csr_waitrequest -> mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_waitrequest
	wire          mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_debugaccess;                          // mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_debugaccess -> dma_subsys:dma_subsys_port8_csr_debugaccess
	wire    [7:0] mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_address;                              // mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_address -> dma_subsys:dma_subsys_port8_csr_address
	wire          mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_read;                                 // mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_read -> dma_subsys:dma_subsys_port8_csr_read
	wire    [3:0] mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_byteenable;                           // mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_byteenable -> dma_subsys:dma_subsys_port8_csr_byteenable
	wire          mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_readdatavalid;                        // dma_subsys:dma_subsys_port8_csr_readdatavalid -> mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_readdatavalid
	wire          mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_write;                                // mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_write -> dma_subsys:dma_subsys_port8_csr_write
	wire   [31:0] mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_writedata;                            // mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_writedata -> dma_subsys:dma_subsys_port8_csr_writedata
	wire    [0:0] mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_burstcount;                           // mm_interconnect_0:dma_subsys_dma_subsys_port8_csr_burstcount -> dma_subsys:dma_subsys_port8_csr_burstcount
	wire  [511:0] mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_readdata;                        // dfd_subsystem:ed_synth_h2f_bridge_s0_readdata -> mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_readdata
	wire          mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_waitrequest;                     // dfd_subsystem:ed_synth_h2f_bridge_s0_waitrequest -> mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_waitrequest
	wire          mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_debugaccess;                     // mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_debugaccess -> dfd_subsystem:ed_synth_h2f_bridge_s0_debugaccess
	wire   [27:0] mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_address;                         // mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_address -> dfd_subsystem:ed_synth_h2f_bridge_s0_address
	wire          mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_read;                            // mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_read -> dfd_subsystem:ed_synth_h2f_bridge_s0_read
	wire   [63:0] mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_byteenable;                      // mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_byteenable -> dfd_subsystem:ed_synth_h2f_bridge_s0_byteenable
	wire          mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_readdatavalid;                   // dfd_subsystem:ed_synth_h2f_bridge_s0_readdatavalid -> mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_readdatavalid
	wire          mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_write;                           // mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_write -> dfd_subsystem:ed_synth_h2f_bridge_s0_write
	wire  [511:0] mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_writedata;                       // mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_writedata -> dfd_subsystem:ed_synth_h2f_bridge_s0_writedata
	wire    [0:0] mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_burstcount;                      // mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_burstcount -> dfd_subsystem:ed_synth_h2f_bridge_s0_burstcount
	wire   [31:0] mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_readdata;                                 // phipps_peak_0:h2f_bridge_s0_readdata -> mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_readdata
	wire          mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_waitrequest;                              // phipps_peak_0:h2f_bridge_s0_waitrequest -> mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_waitrequest
	wire          mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_debugaccess;                              // mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_debugaccess -> phipps_peak_0:h2f_bridge_s0_debugaccess
	wire   [22:0] mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_address;                                  // mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_address -> phipps_peak_0:h2f_bridge_s0_address
	wire          mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_read;                                     // mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_read -> phipps_peak_0:h2f_bridge_s0_read
	wire    [3:0] mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_byteenable;                               // mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_byteenable -> phipps_peak_0:h2f_bridge_s0_byteenable
	wire          mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_readdatavalid;                            // phipps_peak_0:h2f_bridge_s0_readdatavalid -> mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_readdatavalid
	wire          mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_write;                                    // mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_write -> phipps_peak_0:h2f_bridge_s0_write
	wire   [31:0] mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_writedata;                                // mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_writedata -> phipps_peak_0:h2f_bridge_s0_writedata
	wire    [0:0] mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_burstcount;                               // mm_interconnect_0:phipps_peak_0_h2f_bridge_s0_burstcount -> phipps_peak_0:h2f_bridge_s0_burstcount
	wire   [31:0] mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_readdata;             // j204c_f_rx_tx_ip:intel_jesd204c_f_reconfig_xcvr_readdata -> mm_interconnect_0:j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_readdata
	wire          mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_waitrequest;          // j204c_f_rx_tx_ip:intel_jesd204c_f_reconfig_xcvr_waitrequest -> mm_interconnect_0:j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_waitrequest
	wire   [20:0] mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_address;              // mm_interconnect_0:j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_address -> j204c_f_rx_tx_ip:intel_jesd204c_f_reconfig_xcvr_address
	wire          mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_read;                 // mm_interconnect_0:j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_read -> j204c_f_rx_tx_ip:intel_jesd204c_f_reconfig_xcvr_read
	wire    [3:0] mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_byteenable;           // mm_interconnect_0:j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_byteenable -> j204c_f_rx_tx_ip:intel_jesd204c_f_reconfig_xcvr_byteenable
	wire          mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_write;                // mm_interconnect_0:j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_write -> j204c_f_rx_tx_ip:intel_jesd204c_f_reconfig_xcvr_write
	wire   [31:0] mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_writedata;            // mm_interconnect_0:j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_writedata -> j204c_f_rx_tx_ip:intel_jesd204c_f_reconfig_xcvr_writedata
	wire   [31:0] mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_readdata;                           // tod_subsys_0:master_tod_top_0_csr_readdata -> mm_interconnect_0:tod_subsys_0_master_tod_top_0_csr_readdata
	wire          mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_waitrequest;                        // tod_subsys_0:master_tod_top_0_csr_waitrequest -> mm_interconnect_0:tod_subsys_0_master_tod_top_0_csr_waitrequest
	wire    [3:0] mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_address;                            // mm_interconnect_0:tod_subsys_0_master_tod_top_0_csr_address -> tod_subsys_0:master_tod_top_0_csr_address
	wire          mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_read;                               // mm_interconnect_0:tod_subsys_0_master_tod_top_0_csr_read -> tod_subsys_0:master_tod_top_0_csr_read
	wire          mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_write;                              // mm_interconnect_0:tod_subsys_0_master_tod_top_0_csr_write -> tod_subsys_0:master_tod_top_0_csr_write
	wire   [31:0] mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_writedata;                          // mm_interconnect_0:tod_subsys_0_master_tod_top_0_csr_writedata -> tod_subsys_0:master_tod_top_0_csr_writedata
	wire   [31:0] mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_readdata;                 // tod_subsys_0:mtod_subsys_pps_load_tod_0_csr_readdata -> mm_interconnect_0:tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_readdata
	wire          mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_waitrequest;              // tod_subsys_0:mtod_subsys_pps_load_tod_0_csr_waitrequest -> mm_interconnect_0:tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_waitrequest
	wire    [5:0] mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_address;                  // mm_interconnect_0:tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_address -> tod_subsys_0:mtod_subsys_pps_load_tod_0_csr_address
	wire          mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_read;                     // mm_interconnect_0:tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_read -> tod_subsys_0:mtod_subsys_pps_load_tod_0_csr_read
	wire          mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_write;                    // mm_interconnect_0:tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_write -> tod_subsys_0:mtod_subsys_pps_load_tod_0_csr_write
	wire   [31:0] mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_writedata;                // mm_interconnect_0:tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_writedata -> tod_subsys_0:mtod_subsys_pps_load_tod_0_csr_writedata
	wire   [31:0] mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdata;                         // phipps_peak_0:pwr_mtr_h2f_bridge_s0_readdata -> mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdata
	wire          mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_waitrequest;                      // phipps_peak_0:pwr_mtr_h2f_bridge_s0_waitrequest -> mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_waitrequest
	wire          mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_debugaccess;                      // mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_debugaccess -> phipps_peak_0:pwr_mtr_h2f_bridge_s0_debugaccess
	wire   [16:0] mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_address;                          // mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_address -> phipps_peak_0:pwr_mtr_h2f_bridge_s0_address
	wire          mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_read;                             // mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_read -> phipps_peak_0:pwr_mtr_h2f_bridge_s0_read
	wire    [3:0] mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_byteenable;                       // mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_byteenable -> phipps_peak_0:pwr_mtr_h2f_bridge_s0_byteenable
	wire          mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdatavalid;                    // phipps_peak_0:pwr_mtr_h2f_bridge_s0_readdatavalid -> mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdatavalid
	wire          mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_write;                            // mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_write -> phipps_peak_0:pwr_mtr_h2f_bridge_s0_write
	wire   [31:0] mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_writedata;                        // mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_writedata -> phipps_peak_0:pwr_mtr_h2f_bridge_s0_writedata
	wire    [0:0] mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_burstcount;                       // mm_interconnect_0:phipps_peak_0_pwr_mtr_h2f_bridge_s0_burstcount -> phipps_peak_0:pwr_mtr_h2f_bridge_s0_burstcount
	wire          mm_interconnect_0_ftile_debug_status_pio_0_s1_chipselect;                               // mm_interconnect_0:ftile_debug_status_pio_0_s1_chipselect -> ftile_debug_status_pio_0:chipselect
	wire   [31:0] mm_interconnect_0_ftile_debug_status_pio_0_s1_readdata;                                 // ftile_debug_status_pio_0:readdata -> mm_interconnect_0:ftile_debug_status_pio_0_s1_readdata
	wire    [1:0] mm_interconnect_0_ftile_debug_status_pio_0_s1_address;                                  // mm_interconnect_0:ftile_debug_status_pio_0_s1_address -> ftile_debug_status_pio_0:address
	wire          mm_interconnect_0_ftile_debug_status_pio_0_s1_write;                                    // mm_interconnect_0:ftile_debug_status_pio_0_s1_write -> ftile_debug_status_pio_0:write_n
	wire   [31:0] mm_interconnect_0_ftile_debug_status_pio_0_s1_writedata;                                // mm_interconnect_0:ftile_debug_status_pio_0_s1_writedata -> ftile_debug_status_pio_0:writedata
	wire          mm_interconnect_0_ocm_s1_chipselect;                                                    // mm_interconnect_0:ocm_s1_chipselect -> ocm:chipselect
	wire  [127:0] mm_interconnect_0_ocm_s1_readdata;                                                      // ocm:readdata -> mm_interconnect_0:ocm_s1_readdata
	wire   [13:0] mm_interconnect_0_ocm_s1_address;                                                       // mm_interconnect_0:ocm_s1_address -> ocm:address
	wire   [15:0] mm_interconnect_0_ocm_s1_byteenable;                                                    // mm_interconnect_0:ocm_s1_byteenable -> ocm:byteenable
	wire          mm_interconnect_0_ocm_s1_write;                                                         // mm_interconnect_0:ocm_s1_write -> ocm:write
	wire  [127:0] mm_interconnect_0_ocm_s1_writedata;                                                     // mm_interconnect_0:ocm_s1_writedata -> ocm:writedata
	wire          mm_interconnect_0_ocm_s1_clken;                                                         // mm_interconnect_0:ocm_s1_clken -> ocm:clken
	wire          mm_interconnect_0_qsfpdd_status_pio_s1_chipselect;                                      // mm_interconnect_0:qsfpdd_status_pio_s1_chipselect -> qsfpdd_status_pio:chipselect
	wire   [31:0] mm_interconnect_0_qsfpdd_status_pio_s1_readdata;                                        // qsfpdd_status_pio:readdata -> mm_interconnect_0:qsfpdd_status_pio_s1_readdata
	wire    [1:0] mm_interconnect_0_qsfpdd_status_pio_s1_address;                                         // mm_interconnect_0:qsfpdd_status_pio_s1_address -> qsfpdd_status_pio:address
	wire          mm_interconnect_0_qsfpdd_status_pio_s1_write;                                           // mm_interconnect_0:qsfpdd_status_pio_s1_write -> qsfpdd_status_pio:write_n
	wire   [31:0] mm_interconnect_0_qsfpdd_status_pio_s1_writedata;                                       // mm_interconnect_0:qsfpdd_status_pio_s1_writedata -> qsfpdd_status_pio:writedata
	wire          mm_interconnect_0_sys_ctrl_pio_0_s1_chipselect;                                         // mm_interconnect_0:sys_ctrl_pio_0_s1_chipselect -> sys_ctrl_pio_0:chipselect
	wire   [31:0] mm_interconnect_0_sys_ctrl_pio_0_s1_readdata;                                           // sys_ctrl_pio_0:readdata -> mm_interconnect_0:sys_ctrl_pio_0_s1_readdata
	wire    [1:0] mm_interconnect_0_sys_ctrl_pio_0_s1_address;                                            // mm_interconnect_0:sys_ctrl_pio_0_s1_address -> sys_ctrl_pio_0:address
	wire          mm_interconnect_0_sys_ctrl_pio_0_s1_write;                                              // mm_interconnect_0:sys_ctrl_pio_0_s1_write -> sys_ctrl_pio_0:write_n
	wire   [31:0] mm_interconnect_0_sys_ctrl_pio_0_s1_writedata;                                          // mm_interconnect_0:sys_ctrl_pio_0_s1_writedata -> sys_ctrl_pio_0:writedata
	wire    [1:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_awburst;                                       // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awburst -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awburst
	wire    [7:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlen;                                         // hps_sub_sys:agilex_hps_h2f_lw_axi_master_arlen -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlen
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_wstrb;                                         // hps_sub_sys:agilex_hps_h2f_lw_axi_master_wstrb -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_wstrb
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_wready;                                        // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_wready -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_wready
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_rid;                                           // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_rid -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_rid
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_rready;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_rready -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_rready
	wire    [7:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlen;                                         // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awlen -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlen
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_arcache;                                       // hps_sub_sys:agilex_hps_h2f_lw_axi_master_arcache -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arcache
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_wvalid;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_wvalid -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_araddr;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_araddr -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_araddr
	wire    [2:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_arprot;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_arprot -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arprot
	wire    [2:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_awprot;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awprot -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awprot
	wire   [31:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_wdata;                                         // hps_sub_sys:agilex_hps_h2f_lw_axi_master_wdata -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_wdata
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_arvalid;                                       // hps_sub_sys:agilex_hps_h2f_lw_axi_master_arvalid -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_awcache;                                       // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awcache -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awcache
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_arid;                                          // hps_sub_sys:agilex_hps_h2f_lw_axi_master_arid -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arid
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlock;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_arlock -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlock
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlock;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awlock -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlock
	wire   [20:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_awaddr;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awaddr -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_bresp;                                         // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_bresp -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_bresp
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_arready;                                       // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arready -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_arready
	wire   [31:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_rdata;                                         // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_rdata -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_rdata
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_awready;                                       // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awready -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_awready
	wire    [1:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_arburst;                                       // hps_sub_sys:agilex_hps_h2f_lw_axi_master_arburst -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arburst
	wire    [2:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_arsize;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_arsize -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_arsize
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_bready;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_bready -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_bready
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_rlast;                                         // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_rlast -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_rlast
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_wlast;                                         // hps_sub_sys:agilex_hps_h2f_lw_axi_master_wlast -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_wlast
	wire    [1:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_rresp;                                         // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_rresp -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_rresp
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_awid;                                          // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awid -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awid
	wire    [3:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_bid;                                           // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_bid -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_bid
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_bvalid;                                        // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_bvalid -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_bvalid
	wire    [2:0] hps_sub_sys_agilex_hps_h2f_lw_axi_master_awsize;                                        // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awsize -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awsize
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_awvalid;                                       // hps_sub_sys:agilex_hps_h2f_lw_axi_master_awvalid -> mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_awvalid
	wire          hps_sub_sys_agilex_hps_h2f_lw_axi_master_rvalid;                                        // mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_master_rvalid -> hps_sub_sys:agilex_hps_h2f_lw_axi_master_rvalid
	wire   [31:0] jtg_mst_fpga_m_master_readdata;                                                         // mm_interconnect_1:jtg_mst_fpga_m_master_readdata -> jtg_mst:fpga_m_master_readdata
	wire          jtg_mst_fpga_m_master_waitrequest;                                                      // mm_interconnect_1:jtg_mst_fpga_m_master_waitrequest -> jtg_mst:fpga_m_master_waitrequest
	wire   [31:0] jtg_mst_fpga_m_master_address;                                                          // jtg_mst:fpga_m_master_address -> mm_interconnect_1:jtg_mst_fpga_m_master_address
	wire          jtg_mst_fpga_m_master_read;                                                             // jtg_mst:fpga_m_master_read -> mm_interconnect_1:jtg_mst_fpga_m_master_read
	wire    [3:0] jtg_mst_fpga_m_master_byteenable;                                                       // jtg_mst:fpga_m_master_byteenable -> mm_interconnect_1:jtg_mst_fpga_m_master_byteenable
	wire          jtg_mst_fpga_m_master_readdatavalid;                                                    // mm_interconnect_1:jtg_mst_fpga_m_master_readdatavalid -> jtg_mst:fpga_m_master_readdatavalid
	wire          jtg_mst_fpga_m_master_write;                                                            // jtg_mst:fpga_m_master_write -> mm_interconnect_1:jtg_mst_fpga_m_master_write
	wire   [31:0] jtg_mst_fpga_m_master_writedata;                                                        // jtg_mst:fpga_m_master_writedata -> mm_interconnect_1:jtg_mst_fpga_m_master_writedata
	wire   [31:0] mm_interconnect_1_hps_sub_sys_acp_0_csr_readdata;                                       // hps_sub_sys:acp_0_csr_readdata -> mm_interconnect_1:hps_sub_sys_acp_0_csr_readdata
	wire    [0:0] mm_interconnect_1_hps_sub_sys_acp_0_csr_address;                                        // mm_interconnect_1:hps_sub_sys_acp_0_csr_address -> hps_sub_sys:acp_0_csr_address
	wire          mm_interconnect_1_hps_sub_sys_acp_0_csr_read;                                           // mm_interconnect_1:hps_sub_sys_acp_0_csr_read -> hps_sub_sys:acp_0_csr_read
	wire          mm_interconnect_1_hps_sub_sys_acp_0_csr_write;                                          // mm_interconnect_1:hps_sub_sys_acp_0_csr_write -> hps_sub_sys:acp_0_csr_write
	wire   [31:0] mm_interconnect_1_hps_sub_sys_acp_0_csr_writedata;                                      // mm_interconnect_1:hps_sub_sys_acp_0_csr_writedata -> hps_sub_sys:acp_0_csr_writedata
	wire   [31:0] mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_readdata;                              // phipps_peak_0:h2f_lw_bridge_s0_readdata -> mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_readdata
	wire          mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_waitrequest;                           // phipps_peak_0:h2f_lw_bridge_s0_waitrequest -> mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_waitrequest
	wire          mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_debugaccess;                           // mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_debugaccess -> phipps_peak_0:h2f_lw_bridge_s0_debugaccess
	wire   [19:0] mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_address;                               // mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_address -> phipps_peak_0:h2f_lw_bridge_s0_address
	wire          mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_read;                                  // mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_read -> phipps_peak_0:h2f_lw_bridge_s0_read
	wire    [3:0] mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_byteenable;                            // mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_byteenable -> phipps_peak_0:h2f_lw_bridge_s0_byteenable
	wire          mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_readdatavalid;                         // phipps_peak_0:h2f_lw_bridge_s0_readdatavalid -> mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_readdatavalid
	wire          mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_write;                                 // mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_write -> phipps_peak_0:h2f_lw_bridge_s0_write
	wire   [31:0] mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_writedata;                             // mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_writedata -> phipps_peak_0:h2f_lw_bridge_s0_writedata
	wire    [0:0] mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_burstcount;                            // mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_burstcount -> phipps_peak_0:h2f_lw_bridge_s0_burstcount
	wire   [31:0] mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_readdata;                              // dfd_subsystem:h2f_lw_bridge_s0_readdata -> mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_readdata
	wire          mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_waitrequest;                           // dfd_subsystem:h2f_lw_bridge_s0_waitrequest -> mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_waitrequest
	wire          mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_debugaccess;                           // mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_debugaccess -> dfd_subsystem:h2f_lw_bridge_s0_debugaccess
	wire   [12:0] mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_address;                               // mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_address -> dfd_subsystem:h2f_lw_bridge_s0_address
	wire          mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_read;                                  // mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_read -> dfd_subsystem:h2f_lw_bridge_s0_read
	wire    [3:0] mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_byteenable;                            // mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_byteenable -> dfd_subsystem:h2f_lw_bridge_s0_byteenable
	wire          mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_readdatavalid;                         // dfd_subsystem:h2f_lw_bridge_s0_readdatavalid -> mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_readdatavalid
	wire          mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_write;                                 // mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_write -> dfd_subsystem:h2f_lw_bridge_s0_write
	wire   [31:0] mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_writedata;                             // mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_writedata -> dfd_subsystem:h2f_lw_bridge_s0_writedata
	wire    [0:0] mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_burstcount;                            // mm_interconnect_1:dfd_subsystem_h2f_lw_bridge_s0_burstcount -> dfd_subsystem:h2f_lw_bridge_s0_burstcount
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_chipselect;            // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_chipselect -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_rx_avs_chipselect
	wire   [31:0] mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_readdata;              // j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_rx_avs_readdata -> mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_readdata
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_waitrequest;           // j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_rx_avs_waitrequest -> mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_waitrequest
	wire    [9:0] mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_address;               // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_address -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_rx_avs_address
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_read;                  // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_read -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_rx_avs_read
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_write;                 // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_write -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_rx_avs_write
	wire   [31:0] mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_writedata;             // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_writedata -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_rx_avs_writedata
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_chipselect;            // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_chipselect -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_tx_avs_chipselect
	wire   [31:0] mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_readdata;              // j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_tx_avs_readdata -> mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_readdata
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_waitrequest;           // j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_tx_avs_waitrequest -> mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_waitrequest
	wire    [9:0] mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_address;               // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_address -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_tx_avs_address
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_read;                  // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_read -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_tx_avs_read
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_write;                 // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_write -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_tx_avs_write
	wire   [31:0] mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_writedata;             // mm_interconnect_1:j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_writedata -> j204c_f_rx_tx_ip:intel_jesd204c_f_j204c_tx_avs_writedata
	wire   [31:0] mm_interconnect_1_periph_pb_cpu_0_s0_readdata;                                          // periph:pb_cpu_0_s0_readdata -> mm_interconnect_1:periph_pb_cpu_0_s0_readdata
	wire          mm_interconnect_1_periph_pb_cpu_0_s0_waitrequest;                                       // periph:pb_cpu_0_s0_waitrequest -> mm_interconnect_1:periph_pb_cpu_0_s0_waitrequest
	wire          mm_interconnect_1_periph_pb_cpu_0_s0_debugaccess;                                       // mm_interconnect_1:periph_pb_cpu_0_s0_debugaccess -> periph:pb_cpu_0_s0_debugaccess
	wire    [8:0] mm_interconnect_1_periph_pb_cpu_0_s0_address;                                           // mm_interconnect_1:periph_pb_cpu_0_s0_address -> periph:pb_cpu_0_s0_address
	wire          mm_interconnect_1_periph_pb_cpu_0_s0_read;                                              // mm_interconnect_1:periph_pb_cpu_0_s0_read -> periph:pb_cpu_0_s0_read
	wire    [3:0] mm_interconnect_1_periph_pb_cpu_0_s0_byteenable;                                        // mm_interconnect_1:periph_pb_cpu_0_s0_byteenable -> periph:pb_cpu_0_s0_byteenable
	wire          mm_interconnect_1_periph_pb_cpu_0_s0_readdatavalid;                                     // periph:pb_cpu_0_s0_readdatavalid -> mm_interconnect_1:periph_pb_cpu_0_s0_readdatavalid
	wire          mm_interconnect_1_periph_pb_cpu_0_s0_write;                                             // mm_interconnect_1:periph_pb_cpu_0_s0_write -> periph:pb_cpu_0_s0_write
	wire   [31:0] mm_interconnect_1_periph_pb_cpu_0_s0_writedata;                                         // mm_interconnect_1:periph_pb_cpu_0_s0_writedata -> periph:pb_cpu_0_s0_writedata
	wire    [0:0] mm_interconnect_1_periph_pb_cpu_0_s0_burstcount;                                        // mm_interconnect_1:periph_pb_cpu_0_s0_burstcount -> periph:pb_cpu_0_s0_burstcount
	wire   [31:0] mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_readdata;                   // j204c_f_rx_tx_ip:reset_sequencer_0_av_csr_readdata -> mm_interconnect_1:j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_readdata
	wire    [7:0] mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_address;                    // mm_interconnect_1:j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_address -> j204c_f_rx_tx_ip:reset_sequencer_0_av_csr_address
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_read;                       // mm_interconnect_1:j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_read -> j204c_f_rx_tx_ip:reset_sequencer_0_av_csr_read
	wire          mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_write;                      // mm_interconnect_1:j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_write -> j204c_f_rx_tx_ip:reset_sequencer_0_av_csr_write
	wire   [31:0] mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_writedata;                  // mm_interconnect_1:j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_writedata -> j204c_f_rx_tx_ip:reset_sequencer_0_av_csr_writedata
	wire   [31:0] mm_interconnect_1_sys_manager_sysid_control_slave_readdata;                             // sys_manager:sysid_control_slave_readdata -> mm_interconnect_1:sys_manager_sysid_control_slave_readdata
	wire    [0:0] mm_interconnect_1_sys_manager_sysid_control_slave_address;                              // mm_interconnect_1:sys_manager_sysid_control_slave_address -> sys_manager:sysid_control_slave_address
	wire   [31:0] mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata;      // tod_subsys_0:tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata -> mm_interconnect_1:tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata
	wire          mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest;   // tod_subsys_0:tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest -> mm_interconnect_1:tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest
	wire    [4:0] mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_address;       // mm_interconnect_1:tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_address -> tod_subsys_0:tod_timestamp_96b_0_tod_timestamp_96b_csr_address
	wire          mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_read;          // mm_interconnect_1:tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_read -> tod_subsys_0:tod_timestamp_96b_0_tod_timestamp_96b_csr_read
	wire          mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid; // tod_subsys_0:tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid -> mm_interconnect_1:tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid
	wire          mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_write;         // mm_interconnect_1:tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_write -> tod_subsys_0:tod_timestamp_96b_0_tod_timestamp_96b_csr_write
	wire   [31:0] mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata;     // mm_interconnect_1:tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata -> tod_subsys_0:tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata
	wire  [127:0] mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_readdata;                                    // jtg_mst:fpga_m2ocm_pb_s0_readdata -> mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_readdata
	wire          mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_waitrequest;                                 // jtg_mst:fpga_m2ocm_pb_s0_waitrequest -> mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_waitrequest
	wire          mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_debugaccess;                                 // mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_debugaccess -> jtg_mst:fpga_m2ocm_pb_s0_debugaccess
	wire   [17:0] mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_address;                                     // mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_address -> jtg_mst:fpga_m2ocm_pb_s0_address
	wire          mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_read;                                        // mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_read -> jtg_mst:fpga_m2ocm_pb_s0_read
	wire   [15:0] mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_byteenable;                                  // mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_byteenable -> jtg_mst:fpga_m2ocm_pb_s0_byteenable
	wire          mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_readdatavalid;                               // jtg_mst:fpga_m2ocm_pb_s0_readdatavalid -> mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_readdatavalid
	wire          mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_write;                                       // mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_write -> jtg_mst:fpga_m2ocm_pb_s0_write
	wire  [127:0] mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_writedata;                                   // mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_writedata -> jtg_mst:fpga_m2ocm_pb_s0_writedata
	wire    [0:0] mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_burstcount;                                  // mm_interconnect_1:jtg_mst_fpga_m2ocm_pb_s0_burstcount -> jtg_mst:fpga_m2ocm_pb_s0_burstcount
	wire          dma_subsys_dma_ss_master_m0_waitrequest;                                                // mm_interconnect_2:dma_subsys_dma_ss_master_m0_waitrequest -> dma_subsys:dma_ss_master_m0_waitrequest
	wire  [511:0] dma_subsys_dma_ss_master_m0_readdata;                                                   // mm_interconnect_2:dma_subsys_dma_ss_master_m0_readdata -> dma_subsys:dma_ss_master_m0_readdata
	wire          dma_subsys_dma_ss_master_m0_debugaccess;                                                // dma_subsys:dma_ss_master_m0_debugaccess -> mm_interconnect_2:dma_subsys_dma_ss_master_m0_debugaccess
	wire   [36:0] dma_subsys_dma_ss_master_m0_address;                                                    // dma_subsys:dma_ss_master_m0_address -> mm_interconnect_2:dma_subsys_dma_ss_master_m0_address
	wire          dma_subsys_dma_ss_master_m0_read;                                                       // dma_subsys:dma_ss_master_m0_read -> mm_interconnect_2:dma_subsys_dma_ss_master_m0_read
	wire   [63:0] dma_subsys_dma_ss_master_m0_byteenable;                                                 // dma_subsys:dma_ss_master_m0_byteenable -> mm_interconnect_2:dma_subsys_dma_ss_master_m0_byteenable
	wire          dma_subsys_dma_ss_master_m0_readdatavalid;                                              // mm_interconnect_2:dma_subsys_dma_ss_master_m0_readdatavalid -> dma_subsys:dma_ss_master_m0_readdatavalid
	wire    [1:0] dma_subsys_dma_ss_master_m0_response;                                                   // mm_interconnect_2:dma_subsys_dma_ss_master_m0_response -> dma_subsys:dma_ss_master_m0_response
	wire  [511:0] dma_subsys_dma_ss_master_m0_writedata;                                                  // dma_subsys:dma_ss_master_m0_writedata -> mm_interconnect_2:dma_subsys_dma_ss_master_m0_writedata
	wire          dma_subsys_dma_ss_master_m0_write;                                                      // dma_subsys:dma_ss_master_m0_write -> mm_interconnect_2:dma_subsys_dma_ss_master_m0_write
	wire          dma_subsys_dma_ss_master_m0_writeresponsevalid;                                         // mm_interconnect_2:dma_subsys_dma_ss_master_m0_writeresponsevalid -> dma_subsys:dma_ss_master_m0_writeresponsevalid
	wire    [4:0] dma_subsys_dma_ss_master_m0_burstcount;                                                 // dma_subsys:dma_ss_master_m0_burstcount -> mm_interconnect_2:dma_subsys_dma_ss_master_m0_burstcount
	wire          dma_subsys_ext_hps_m_master_expanded_master_waitrequest;                                // mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_waitrequest -> dma_subsys:ext_hps_m_master_expanded_master_waitrequest
	wire   [31:0] dma_subsys_ext_hps_m_master_expanded_master_readdata;                                   // mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_readdata -> dma_subsys:ext_hps_m_master_expanded_master_readdata
	wire   [36:0] dma_subsys_ext_hps_m_master_expanded_master_address;                                    // dma_subsys:ext_hps_m_master_expanded_master_address -> mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_address
	wire          dma_subsys_ext_hps_m_master_expanded_master_read;                                       // dma_subsys:ext_hps_m_master_expanded_master_read -> mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_read
	wire    [3:0] dma_subsys_ext_hps_m_master_expanded_master_byteenable;                                 // dma_subsys:ext_hps_m_master_expanded_master_byteenable -> mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_byteenable
	wire          dma_subsys_ext_hps_m_master_expanded_master_readdatavalid;                              // mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_readdatavalid -> dma_subsys:ext_hps_m_master_expanded_master_readdatavalid
	wire          dma_subsys_ext_hps_m_master_expanded_master_write;                                      // dma_subsys:ext_hps_m_master_expanded_master_write -> mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_write
	wire   [31:0] dma_subsys_ext_hps_m_master_expanded_master_writedata;                                  // dma_subsys:ext_hps_m_master_expanded_master_writedata -> mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_writedata
	wire    [0:0] dma_subsys_ext_hps_m_master_expanded_master_burstcount;                                 // dma_subsys:ext_hps_m_master_expanded_master_burstcount -> mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_burstcount
	wire    [1:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_awburst;                                         // mm_interconnect_2:hps_sub_sys_acp_0_s0_awburst -> hps_sub_sys:acp_0_s0_awburst
	wire    [7:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_arlen;                                           // mm_interconnect_2:hps_sub_sys_acp_0_s0_arlen -> hps_sub_sys:acp_0_s0_arlen
	wire   [63:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_wstrb;                                           // mm_interconnect_2:hps_sub_sys_acp_0_s0_wstrb -> hps_sub_sys:acp_0_s0_wstrb
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_wready;                                          // hps_sub_sys:acp_0_s0_wready -> mm_interconnect_2:hps_sub_sys_acp_0_s0_wready
	wire    [3:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_rid;                                             // hps_sub_sys:acp_0_s0_rid -> mm_interconnect_2:hps_sub_sys_acp_0_s0_rid
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_rready;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_rready -> hps_sub_sys:acp_0_s0_rready
	wire    [7:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_awlen;                                           // mm_interconnect_2:hps_sub_sys_acp_0_s0_awlen -> hps_sub_sys:acp_0_s0_awlen
	wire    [3:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_arcache;                                         // mm_interconnect_2:hps_sub_sys_acp_0_s0_arcache -> hps_sub_sys:acp_0_s0_arcache
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_wvalid;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_wvalid -> hps_sub_sys:acp_0_s0_wvalid
	wire   [36:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_araddr;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_araddr -> hps_sub_sys:acp_0_s0_araddr
	wire    [2:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_arprot;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_arprot -> hps_sub_sys:acp_0_s0_arprot
	wire    [2:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_awprot;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_awprot -> hps_sub_sys:acp_0_s0_awprot
	wire  [511:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_wdata;                                           // mm_interconnect_2:hps_sub_sys_acp_0_s0_wdata -> hps_sub_sys:acp_0_s0_wdata
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_arvalid;                                         // mm_interconnect_2:hps_sub_sys_acp_0_s0_arvalid -> hps_sub_sys:acp_0_s0_arvalid
	wire    [3:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_awcache;                                         // mm_interconnect_2:hps_sub_sys_acp_0_s0_awcache -> hps_sub_sys:acp_0_s0_awcache
	wire    [3:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_arid;                                            // mm_interconnect_2:hps_sub_sys_acp_0_s0_arid -> hps_sub_sys:acp_0_s0_arid
	wire    [0:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_arlock;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_arlock -> hps_sub_sys:acp_0_s0_arlock
	wire    [0:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_awlock;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_awlock -> hps_sub_sys:acp_0_s0_awlock
	wire   [36:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_awaddr;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_awaddr -> hps_sub_sys:acp_0_s0_awaddr
	wire    [1:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_bresp;                                           // hps_sub_sys:acp_0_s0_bresp -> mm_interconnect_2:hps_sub_sys_acp_0_s0_bresp
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_arready;                                         // hps_sub_sys:acp_0_s0_arready -> mm_interconnect_2:hps_sub_sys_acp_0_s0_arready
	wire  [511:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_rdata;                                           // hps_sub_sys:acp_0_s0_rdata -> mm_interconnect_2:hps_sub_sys_acp_0_s0_rdata
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_awready;                                         // hps_sub_sys:acp_0_s0_awready -> mm_interconnect_2:hps_sub_sys_acp_0_s0_awready
	wire    [1:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_arburst;                                         // mm_interconnect_2:hps_sub_sys_acp_0_s0_arburst -> hps_sub_sys:acp_0_s0_arburst
	wire    [2:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_arsize;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_arsize -> hps_sub_sys:acp_0_s0_arsize
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_bready;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_bready -> hps_sub_sys:acp_0_s0_bready
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_rlast;                                           // hps_sub_sys:acp_0_s0_rlast -> mm_interconnect_2:hps_sub_sys_acp_0_s0_rlast
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_wlast;                                           // mm_interconnect_2:hps_sub_sys_acp_0_s0_wlast -> hps_sub_sys:acp_0_s0_wlast
	wire    [1:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_rresp;                                           // hps_sub_sys:acp_0_s0_rresp -> mm_interconnect_2:hps_sub_sys_acp_0_s0_rresp
	wire    [3:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_awid;                                            // mm_interconnect_2:hps_sub_sys_acp_0_s0_awid -> hps_sub_sys:acp_0_s0_awid
	wire    [3:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_bid;                                             // hps_sub_sys:acp_0_s0_bid -> mm_interconnect_2:hps_sub_sys_acp_0_s0_bid
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_bvalid;                                          // hps_sub_sys:acp_0_s0_bvalid -> mm_interconnect_2:hps_sub_sys_acp_0_s0_bvalid
	wire    [2:0] mm_interconnect_2_hps_sub_sys_acp_0_s0_awsize;                                          // mm_interconnect_2:hps_sub_sys_acp_0_s0_awsize -> hps_sub_sys:acp_0_s0_awsize
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_awvalid;                                         // mm_interconnect_2:hps_sub_sys_acp_0_s0_awvalid -> hps_sub_sys:acp_0_s0_awvalid
	wire          mm_interconnect_2_hps_sub_sys_acp_0_s0_rvalid;                                          // hps_sub_sys:acp_0_s0_rvalid -> mm_interconnect_2:hps_sub_sys_acp_0_s0_rvalid
	wire   [31:0] jtg_mst_hps_m_master_readdata;                                                          // mm_interconnect_3:jtg_mst_hps_m_master_readdata -> jtg_mst:hps_m_master_readdata
	wire          jtg_mst_hps_m_master_waitrequest;                                                       // mm_interconnect_3:jtg_mst_hps_m_master_waitrequest -> jtg_mst:hps_m_master_waitrequest
	wire   [31:0] jtg_mst_hps_m_master_address;                                                           // jtg_mst:hps_m_master_address -> mm_interconnect_3:jtg_mst_hps_m_master_address
	wire          jtg_mst_hps_m_master_read;                                                              // jtg_mst:hps_m_master_read -> mm_interconnect_3:jtg_mst_hps_m_master_read
	wire    [3:0] jtg_mst_hps_m_master_byteenable;                                                        // jtg_mst:hps_m_master_byteenable -> mm_interconnect_3:jtg_mst_hps_m_master_byteenable
	wire          jtg_mst_hps_m_master_readdatavalid;                                                     // mm_interconnect_3:jtg_mst_hps_m_master_readdatavalid -> jtg_mst:hps_m_master_readdatavalid
	wire          jtg_mst_hps_m_master_write;                                                             // jtg_mst:hps_m_master_write -> mm_interconnect_3:jtg_mst_hps_m_master_write
	wire   [31:0] jtg_mst_hps_m_master_writedata;                                                         // jtg_mst:hps_m_master_writedata -> mm_interconnect_3:jtg_mst_hps_m_master_writedata
	wire   [31:0] mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_readdata;                  // dma_subsys:ext_hps_m_master_windowed_slave_readdata -> mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_readdata
	wire          mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_waitrequest;               // dma_subsys:ext_hps_m_master_windowed_slave_waitrequest -> mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_waitrequest
	wire   [29:0] mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_address;                   // mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_address -> dma_subsys:ext_hps_m_master_windowed_slave_address
	wire          mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_read;                      // mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_read -> dma_subsys:ext_hps_m_master_windowed_slave_read
	wire    [3:0] mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_byteenable;                // mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_byteenable -> dma_subsys:ext_hps_m_master_windowed_slave_byteenable
	wire          mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_readdatavalid;             // dma_subsys:ext_hps_m_master_windowed_slave_readdatavalid -> mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_readdatavalid
	wire          mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_write;                     // mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_write -> dma_subsys:ext_hps_m_master_windowed_slave_write
	wire   [31:0] mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_writedata;                 // mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_writedata -> dma_subsys:ext_hps_m_master_windowed_slave_writedata
	wire    [0:0] mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_burstcount;                // mm_interconnect_3:dma_subsys_ext_hps_m_master_windowed_slave_burstcount -> dma_subsys:ext_hps_m_master_windowed_slave_burstcount
	wire          irq_mapper_receiver2_irq;                                                               // dma_subsys:dma_subsys_port8_rx_dma_ch1_irq_irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                               // dma_subsys:dma_subsys_port8_tx_dma_ch1_irq_irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                               // phipps_peak_0:fifo_full_intr_irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                               // ftile_debug_status_pio_0:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                               // qsfpdd_status_pio:irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                                               // phipps_peak_0:lphy_ss_top_0_lphy_ss_top_pwr_mtr_fft_hist_done_intr_l1_irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                                               // phipps_peak_0:lphy_ss_top_0_lphy_ss_top_pwr_mtr_fft_hist_done_intr_l2_irq -> irq_mapper:receiver8_irq
	wire          irq_mapper_receiver9_irq;                                                               // phipps_peak_0:lphy_ss_top_0_lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l1_irq -> irq_mapper:receiver9_irq
	wire          irq_mapper_receiver10_irq;                                                              // phipps_peak_0:lphy_ss_top_0_lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l2_irq -> irq_mapper:receiver10_irq
	wire          irq_mapper_receiver11_irq;                                                              // tod_subsys_0:mtod_subsys_pps_load_tod_0_pps_irq_irq -> irq_mapper:receiver11_irq
	wire          irq_mapper_receiver12_irq;                                                              // phipps_peak_0:timeout_cntr_intr_cplane_irq -> irq_mapper:receiver12_irq
	wire          irq_mapper_receiver13_irq;                                                              // phipps_peak_0:timeout_cntr_intr_uplane_irq -> irq_mapper:receiver13_irq
	wire   [31:0] hps_sub_sys_agilex_hps_f2h_irq0_irq;                                                    // irq_mapper:sender_irq -> hps_sub_sys:agilex_hps_f2h_irq0_irq
	wire    [1:0] periph_ilc_irq_irq;                                                                     // irq_mapper_001:sender_irq -> periph:ILC_irq_irq
	wire          irq_mapper_receiver0_irq;                                                               // periph:button_pio_irq_irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire          irq_mapper_receiver1_irq;                                                               // periph:dipsw_pio_irq_irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	wire          rst_controller_reset_out_reset;                                                         // rst_controller:reset_out -> [dma_subsys:dma_rst_100_in_reset_reset, ftile_debug_status_pio_0:reset_n, hps_sub_sys:acp_0_csr_reset_reset, hps_sub_sys:agilex_hps_h2f_axi_reset_reset_n, hps_sub_sys:agilex_hps_h2f_lw_axi_reset_reset_n, hssi_ss_1:app_ss_lite_areset_n, irq_mapper_001:reset, j204c_f_rx_tx_ip:mgmt_reset_in_reset_reset_n, ocm:reset, qsfpdd_status_pio:reset_n, rst_translator:in_reset, sys_ctrl_pio_0:reset_n, sys_manager:sysid_reset_reset_n, tod_subsys_0:mtod_subsys_rstn_in_reset_reset_n]
	wire          rst_controller_reset_out_reset_req;                                                     // rst_controller:reset_req -> [ocm:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                                     // rst_controller_001:reset_out -> hps_sub_sys:acp_0_reset_reset
	wire          rst_controller_002_reset_out_reset;                                                     // rst_controller_002:reset_out -> [jtg_mst:reset_reset_n, mm_interconnect_0:hps_sub_sys_agilex_hps_h2f_axi_reset_reset_bridge_in_reset_reset, mm_interconnect_0:jtg_mst_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_sub_sys_agilex_hps_h2f_lw_axi_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtg_mst_reset_reset_bridge_in_reset_reset, mm_interconnect_2:crosser_002_in_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:dma_subsys_ext_hps_m_master_expanded_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:jtg_mst_reset_reset_bridge_in_reset_reset, periph:reset_reset_n, tod_subsys_0:master_tod_top_0_i_reconfig_rst_n_reset_n, tod_subsys_0:tod_slave_tod_subsys_rst_100_in_reset_reset_n]
	wire          rst_controller_003_reset_out_reset;                                                     // rst_controller_003:reset_out -> rst_ss_0:reset_bridge_rec_rx_in_reset_reset
	wire          rst_controller_004_reset_out_reset;                                                     // rst_controller_004:reset_out -> rst_ss_0:reset_bridge_tx_div_in_reset_reset
	wire          rst_controller_005_reset_out_reset;                                                     // rst_controller_005:reset_out -> [tod_subsys_0:mtod_subsys_pps_load_tod_0_csr_reset_reset, tod_subsys_0:mtod_subsys_pps_load_tod_0_reset_reset, tod_subsys_0:reset_bridge_156_in_reset_reset]
	wire          rst_controller_006_reset_out_reset;                                                     // rst_controller_006:reset_out -> [mm_interconnect_0:dfd_subsystem_ed_synth_h2f_bridge_s0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:dfd_subsystem_reset_csr_reset_bridge_in_reset_reset, mm_interconnect_1:phipps_peak_0_csr_in_reset_reset_bridge_in_reset_reset, mm_interconnect_1:phipps_peak_0_h2f_lw_bridge_s0_translator_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_007_reset_out_reset;                                                     // rst_controller_007:reset_out -> [mm_interconnect_2:dma_subsys_dma_rst_100_in_reset_reset_bridge_in_reset_reset, mm_interconnect_2:dma_subsys_dma_ss_master_m0_translator_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_008_reset_out_reset;                                                     // rst_controller_008:reset_out -> [mm_interconnect_2:hps_sub_sys_acp_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_sub_sys_acp_0_s0_translator_clk_reset_reset_bridge_in_reset_reset]

	ftile_debug_status_pio_0 ftile_debug_status_pio_0 (
		.clk        (sys_manager_clk_100_out_clk_clk),                          //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_0_ftile_debug_status_pio_0_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_0_ftile_debug_status_pio_0_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_0_ftile_debug_status_pio_0_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_0_ftile_debug_status_pio_0_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_0_ftile_debug_status_pio_0_s1_readdata),   //  output,  width = 32,                    .readdata
		.in_port    (ftile_debug_status_econ_export),                           //   input,  width = 20, external_connection.export
		.irq        (irq_mapper_receiver5_irq)                                  //  output,   width = 1,                 irq.irq
	);

	hssi_ss_1 hssi_ss_1 (
		.app_ss_lite_clk                    (sys_manager_clk_100_out_clk_clk),                                  //   input,    width = 1,                         axi4_lite_clk.clk
		.app_ss_lite_areset_n               (~rst_controller_reset_out_reset),                                  //   input,    width = 1,                       axi4_lite_reset.reset_n
		.app_ss_lite_awaddr                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awaddr),           //   input,   width = 26,                   axi4_lite_interface.awaddr
		.app_ss_lite_awprot                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awprot),           //   input,    width = 3,                                      .awprot
		.app_ss_lite_awvalid                (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awvalid),          //   input,    width = 1,                                      .awvalid
		.ss_app_lite_awready                (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awready),          //  output,    width = 1,                                      .awready
		.app_ss_lite_wdata                  (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wdata),            //   input,   width = 32,                                      .wdata
		.app_ss_lite_wstrb                  (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wstrb),            //   input,    width = 4,                                      .wstrb
		.app_ss_lite_wvalid                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wvalid),           //   input,    width = 1,                                      .wvalid
		.ss_app_lite_wready                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wready),           //  output,    width = 1,                                      .wready
		.ss_app_lite_bresp                  (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bresp),            //  output,    width = 2,                                      .bresp
		.ss_app_lite_bvalid                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bvalid),           //  output,    width = 1,                                      .bvalid
		.app_ss_lite_bready                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bready),           //   input,    width = 1,                                      .bready
		.app_ss_lite_araddr                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_araddr),           //   input,   width = 26,                                      .araddr
		.app_ss_lite_arprot                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arprot),           //   input,    width = 3,                                      .arprot
		.app_ss_lite_arvalid                (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arvalid),          //   input,    width = 1,                                      .arvalid
		.ss_app_lite_arready                (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arready),          //  output,    width = 1,                                      .arready
		.ss_app_lite_rdata                  (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rdata),            //  output,   width = 32,                                      .rdata
		.ss_app_lite_rvalid                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rvalid),           //  output,    width = 1,                                      .rvalid
		.app_ss_lite_rready                 (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rready),           //   input,    width = 1,                                      .rready
		.ss_app_lite_rresp                  (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rresp),            //  output,    width = 2,                                      .rresp
		.p0_app_ss_st_tx_clk                (clk_ss_0_clk_ftile_402_out_clk_clk),                               //   input,    width = 1,                      p0_axi_st_tx_clk.clk
		.p0_app_ss_st_tx_areset_n           (hssi_ss_1_p0_axi_st_tx_reset_reset_n),                             //   input,    width = 1,                    p0_axi_st_tx_reset.reset_n
		.p0_app_ss_st_tx_tvalid             (hssi_ss_1_p0_axi_st_tx_interface_tvalid),                          //   input,    width = 1,                p0_axi_st_tx_interface.tvalid
		.p0_ss_app_st_tx_tready             (hssi_ss_1_p0_axi_st_tx_interface_tready),                          //  output,    width = 1,                                      .tready
		.p0_app_ss_st_tx_tdata              (hssi_ss_1_p0_axi_st_tx_interface_tdata),                           //   input,   width = 64,                                      .tdata
		.p0_app_ss_st_tx_tkeep              (hssi_ss_1_p0_axi_st_tx_interface_tkeep),                           //   input,    width = 8,                                      .tkeep
		.p0_app_ss_st_tx_tlast              (hssi_ss_1_p0_axi_st_tx_interface_tlast),                           //   input,    width = 1,                                      .tlast
		.p0_app_ss_st_tx_tuser_client       (hssi_ss_1_p0_axi_st_tx_interface_tuser),                           //   input,    width = 2,                                      .tuser
		.p0_app_ss_st_tx_tuser_ptp          (hssi_ss_1_p0_tx_tuser_ptp_tuser_1),                                //   input,   width = 94,                       p0_tx_tuser_ptp.tuser_1
		.p0_app_ss_st_tx_tuser_ptp_extended (hssi_ss_1_p0_tx_tuser_ptp_extended_tuser_2),                       //   input,  width = 328,              p0_tx_tuser_ptp_extended.tuser_2
		.p0_app_ss_st_tx_tuser_last_segment (hssi_ss_1_p0_axi_st_tx_tuser_last_seg_interface_tx_last_segment),  //   input,    width = 1, p0_axi_st_tx_tuser_last_seg_interface.tx_last_segment
		.p0_app_ss_st_rx_clk                (clk_ss_0_clk_ftile_402_out_clk_clk),                               //   input,    width = 1,                      p0_axi_st_rx_clk.clk
		.p0_app_ss_st_rx_areset_n           (hssi_ss_1_p0_axi_st_rx_reset_reset_n),                             //   input,    width = 1,                    p0_axi_st_rx_reset.reset_n
		.p0_ss_app_st_rx_tvalid             (hssi_ss_1_p0_axi_st_rx_interface_tvalid),                          //  output,    width = 1,                p0_axi_st_rx_interface.tvalid
		.p0_ss_app_st_rx_tdata              (hssi_ss_1_p0_axi_st_rx_interface_tdata),                           //  output,   width = 64,                                      .tdata
		.p0_ss_app_st_rx_tkeep              (hssi_ss_1_p0_axi_st_rx_interface_tkeep),                           //  output,    width = 8,                                      .tkeep
		.p0_ss_app_st_rx_tlast              (hssi_ss_1_p0_axi_st_rx_interface_tlast),                           //  output,    width = 1,                                      .tlast
		.p0_ss_app_st_rx_tuser_client       (hssi_ss_1_p0_axi_st_rx_interface_tuser),                           //  output,    width = 7,                                      .tuser
		.p0_ss_app_st_rx_tuser_last_segment (),                                                                 //  output,    width = 1, p0_axi_st_rx_tuser_last_seg_interface.rx_last_segment
		.p0_ss_app_st_rx_tuser_sts          (hssi_ss_1_p0_rx_tuser_status_tuser_1),                             //  output,    width = 5,                    p0_rx_tuser_status.tuser_1
		.p0_app_ss_st_txtod_tvalid          (tod_subsys_0_tod_slave_port_8_tod_stack_tx_tod_interface_tvalid),  //   input,    width = 1,            p0_axi_st_tx_ptp_interface.tvalid
		.p0_app_ss_st_txtod_tdata           (tod_subsys_0_tod_slave_port_8_tod_stack_tx_tod_interface_tdata),   //   input,   width = 96,                                      .tdata
		.p0_app_ss_st_rxtod_tvalid          (tod_subsys_0_tod_slave_port_8_tod_stack_rx_tod_interface_tvalid),  //   input,    width = 1,            p0_axi_st_rx_ptp_interface.tvalid
		.p0_app_ss_st_rxtod_tdata           (tod_subsys_0_tod_slave_port_8_tod_stack_rx_tod_interface_tdata),   //   input,   width = 96,                                      .tdata
		.p0_ss_app_st_txegrts0_tvalid       (hssi_ss_1_p0_axi_st_tx_egrs0_interface_tvalid),                    //  output,    width = 1,          p0_axi_st_tx_egrs0_interface.tvalid
		.p0_ss_app_st_txegrts0_tdata        (hssi_ss_1_p0_axi_st_tx_egrs0_interface_tdata),                     //  output,  width = 128,                                      .tdata
		.p0_ss_app_st_rxingrts0_tvalid      (hssi_ss_1_p0_axi_st_rx_ingrs0_interface_tvalid),                   //  output,    width = 1,         p0_axi_st_rx_ingrs0_interface.tvalid
		.p0_ss_app_st_rxingrts0_tdata       (hssi_ss_1_p0_axi_st_rx_ingrs0_interface_tdata),                    //  output,   width = 96,                                      .tdata
		.i_p0_tx_pause                      (hssi_ss_1_p0_tx_flow_control_interface_i_p0_tx_pause),             //   input,    width = 1,          p0_tx_flow_control_interface.i_p0_tx_pause
		.i_p0_tx_pfc                        (hssi_ss_1_p0_tx_flow_control_interface_i_p0_tx_pfc),               //   input,    width = 8,                                      .i_p0_tx_pfc
		.o_p0_rx_pause                      (),                                                                 //  output,    width = 1,          p0_rx_flow_control_interface.o_p0_rx_pause
		.o_p0_rx_pfc                        (),                                                                 //  output,    width = 8,                                      .o_p0_rx_pfc
		.p0_tx_serial                       (hssi_ss_1_p0_tx_srl_interface_p0_tx_serial),                       //  output,    width = 1,                   p0_tx_srl_interface.p0_tx_serial
		.p0_tx_serial_n                     (hssi_ss_1_p0_tx_srl_interface_p0_tx_serial_n),                     //  output,    width = 1,                                      .p0_tx_serial_n
		.p0_rx_serial                       (hssi_ss_1_p0_rx_srl_interface_p0_rx_serial),                       //   input,    width = 1,                   p0_rx_srl_interface.p0_rx_serial
		.p0_rx_serial_n                     (hssi_ss_1_p0_rx_srl_interface_p0_rx_serial_n),                     //   input,    width = 1,                                      .p0_rx_serial_n
		.port0_led_speed                    (hssi_ss_1_p0_qsfp_led_sts_if_port0_led_speed),                     //  output,    width = 3,                    p0_qsfp_led_sts_if.port0_led_speed
		.port0_led_status                   (hssi_ss_1_p0_qsfp_led_sts_if_port0_led_status),                    //  output,    width = 3,                                      .port0_led_status
		.port1_led_speed                    (hssi_ss_1_p1_qsfp_led_sts_if_port1_led_speed),                     //  output,    width = 3,                    p1_qsfp_led_sts_if.port1_led_speed
		.port1_led_status                   (hssi_ss_1_p1_qsfp_led_sts_if_port1_led_status),                    //  output,    width = 3,                                      .port1_led_status
		.port2_led_speed                    (hssi_ss_1_p2_qsfp_led_sts_if_port2_led_speed),                     //  output,    width = 3,                    p2_qsfp_led_sts_if.port2_led_speed
		.port2_led_status                   (hssi_ss_1_p2_qsfp_led_sts_if_port2_led_status),                    //  output,    width = 3,                                      .port2_led_status
		.port3_led_speed                    (hssi_ss_1_p3_qsfp_led_sts_if_port3_led_speed),                     //  output,    width = 3,                    p3_qsfp_led_sts_if.port3_led_speed
		.port3_led_status                   (hssi_ss_1_p3_qsfp_led_sts_if_port3_led_status),                    //  output,    width = 3,                                      .port3_led_status
		.port4_led_speed                    (hssi_ss_1_p4_qsfp_led_sts_if_port4_led_speed),                     //  output,    width = 3,                    p4_qsfp_led_sts_if.port4_led_speed
		.port4_led_status                   (hssi_ss_1_p4_qsfp_led_sts_if_port4_led_status),                    //  output,    width = 3,                                      .port4_led_status
		.port5_led_speed                    (hssi_ss_1_p5_qsfp_led_sts_if_port5_led_speed),                     //  output,    width = 3,                    p5_qsfp_led_sts_if.port5_led_speed
		.port5_led_status                   (hssi_ss_1_p5_qsfp_led_sts_if_port5_led_status),                    //  output,    width = 3,                                      .port5_led_status
		.port6_led_speed                    (hssi_ss_1_p6_qsfp_led_sts_if_port6_led_speed),                     //  output,    width = 3,                    p6_qsfp_led_sts_if.port6_led_speed
		.port6_led_status                   (hssi_ss_1_p6_qsfp_led_sts_if_port6_led_status),                    //  output,    width = 3,                                      .port6_led_status
		.port7_led_speed                    (hssi_ss_1_p7_qsfp_led_sts_if_port7_led_speed),                     //  output,    width = 3,                    p7_qsfp_led_sts_if.port7_led_speed
		.port7_led_status                   (hssi_ss_1_p7_qsfp_led_sts_if_port7_led_status),                    //  output,    width = 3,                                      .port7_led_status
		.port8_led_speed                    (hssi_ss_1_p8_qsfp_led_sts_if_port8_led_speed),                     //  output,    width = 3,                    p8_qsfp_led_sts_if.port8_led_speed
		.port8_led_status                   (hssi_ss_1_p8_qsfp_led_sts_if_port8_led_status),                    //  output,    width = 3,                                      .port8_led_status
		.port9_led_speed                    (hssi_ss_1_p9_qsfp_led_sts_if_port9_led_speed),                     //  output,    width = 3,                    p9_qsfp_led_sts_if.port9_led_speed
		.port9_led_status                   (hssi_ss_1_p9_qsfp_led_sts_if_port9_led_status),                    //  output,    width = 3,                                      .port9_led_status
		.port10_led_speed                   (hssi_ss_1_p10_qsfp_led_sts_if_port10_led_speed),                   //  output,    width = 3,                   p10_qsfp_led_sts_if.port10_led_speed
		.port10_led_status                  (hssi_ss_1_p10_qsfp_led_sts_if_port10_led_status),                  //  output,    width = 3,                                      .port10_led_status
		.port11_led_speed                   (hssi_ss_1_p11_qsfp_led_sts_if_port11_led_speed),                   //  output,    width = 3,                   p11_qsfp_led_sts_if.port11_led_speed
		.port11_led_status                  (hssi_ss_1_p11_qsfp_led_sts_if_port11_led_status),                  //  output,    width = 3,                                      .port11_led_status
		.port12_led_speed                   (hssi_ss_1_p12_qsfp_led_sts_if_port12_led_speed),                   //  output,    width = 3,                   p12_qsfp_led_sts_if.port12_led_speed
		.port12_led_status                  (hssi_ss_1_p12_qsfp_led_sts_if_port12_led_status),                  //  output,    width = 3,                                      .port12_led_status
		.port13_led_speed                   (hssi_ss_1_p13_qsfp_led_sts_if_port13_led_speed),                   //  output,    width = 3,                   p13_qsfp_led_sts_if.port13_led_speed
		.port13_led_status                  (hssi_ss_1_p13_qsfp_led_sts_if_port13_led_status),                  //  output,    width = 3,                                      .port13_led_status
		.port14_led_speed                   (hssi_ss_1_p14_qsfp_led_sts_if_port14_led_speed),                   //  output,    width = 3,                   p14_qsfp_led_sts_if.port14_led_speed
		.port14_led_status                  (hssi_ss_1_p14_qsfp_led_sts_if_port14_led_status),                  //  output,    width = 3,                                      .port14_led_status
		.port15_led_speed                   (hssi_ss_1_p15_qsfp_led_sts_if_port15_led_speed),                   //  output,    width = 3,                   p15_qsfp_led_sts_if.port15_led_speed
		.port15_led_status                  (hssi_ss_1_p15_qsfp_led_sts_if_port15_led_status),                  //  output,    width = 3,                                      .port15_led_status
		.port16_led_speed                   (hssi_ss_1_p16_qsfp_led_sts_if_port16_led_speed),                   //  output,    width = 3,                   p16_qsfp_led_sts_if.port16_led_speed
		.port16_led_status                  (hssi_ss_1_p16_qsfp_led_sts_if_port16_led_status),                  //  output,    width = 3,                                      .port16_led_status
		.port17_led_speed                   (hssi_ss_1_p17_qsfp_led_sts_if_port17_led_speed),                   //  output,    width = 3,                   p17_qsfp_led_sts_if.port17_led_speed
		.port17_led_status                  (hssi_ss_1_p17_qsfp_led_sts_if_port17_led_status),                  //  output,    width = 3,                                      .port17_led_status
		.port18_led_speed                   (hssi_ss_1_p18_qsfp_led_sts_if_port18_led_speed),                   //  output,    width = 3,                   p18_qsfp_led_sts_if.port18_led_speed
		.port18_led_status                  (hssi_ss_1_p18_qsfp_led_sts_if_port18_led_status),                  //  output,    width = 3,                                      .port18_led_status
		.port19_led_speed                   (hssi_ss_1_p19_qsfp_led_sts_if_port19_led_speed),                   //  output,    width = 3,                   p19_qsfp_led_sts_if.port19_led_speed
		.port19_led_status                  (hssi_ss_1_p19_qsfp_led_sts_if_port19_led_status),                  //  output,    width = 3,                                      .port19_led_status
		.p0_tx_lanes_stable                 (hssi_ss_1_p0_misc_interface_p0_tx_lanes_stable),                   //  output,    width = 1,                     p0_misc_interface.p0_tx_lanes_stable
		.p0_rx_pcs_ready                    (hssi_ss_1_p0_misc_interface_p0_rx_pcs_ready),                      //  output,    width = 1,                                      .p0_rx_pcs_ready
		.o_p0_tx_pll_locked                 (hssi_ss_1_p0_misc_interface_o_p0_tx_pll_locked),                   //  output,    width = 1,                                      .o_p0_tx_pll_locked
		.o_p0_rx_pcs_fully_aligned          (),                                                                 //  output,    width = 1,               p0_rx_pcs_fully_aligned.o_p0_rx_pcs_fully_aligned
		.o_p0_tx_ptp_ready                  (hssi_ss_1_p0_tx_ptp_ready_o_p0_tx_ptp_ready),                      //  output,    width = 1,                       p0_tx_ptp_ready.o_p0_tx_ptp_ready
		.o_p0_rx_ptp_ready                  (hssi_ss_1_p0_rx_ptp_ready_o_p0_rx_ptp_ready),                      //  output,    width = 1,                       p0_rx_ptp_ready.o_p0_rx_ptp_ready
		.o_p0_rx_ptp_offset_data_valid      (hssi_ss_1_p0_ptp_offset_data_valid_o_p0_rx_ptp_offset_data_valid), //  output,    width = 1,              p0_ptp_offset_data_valid.o_p0_rx_ptp_offset_data_valid
		.o_p0_tx_ptp_offset_data_valid      (hssi_ss_1_p0_ptp_offset_data_valid_o_p0_tx_ptp_offset_data_valid), //  output,    width = 1,                                      .o_p0_tx_ptp_offset_data_valid
		.subsystem_cold_rst_n               (hssi_ss_1_subsystem_cold_rst_n_reset_n),                           //   input,    width = 1,                  subsystem_cold_rst_n.reset_n
		.subsystem_cold_rst_ack_n           (hssi_ss_1_subsystem_cold_rst_ack_n_reset_n),                       //  output,    width = 1,              subsystem_cold_rst_ack_n.reset_n
		.i_p0_tx_rst_n                      (hssi_ss_1_i_p0_tx_rst_n_reset_n),                                  //   input,    width = 1,                         i_p0_tx_rst_n.reset_n
		.i_p0_rx_rst_n                      (hssi_ss_1_i_p0_rx_rst_n_reset_n),                                  //   input,    width = 1,                         i_p0_rx_rst_n.reset_n
		.o_p0_rx_rst_ack_n                  (hssi_ss_1_o_p0_rx_rst_ack_n_reset_n),                              //  output,    width = 1,                     o_p0_rx_rst_ack_n.reset_n
		.o_p0_tx_rst_ack_n                  (hssi_ss_1_o_p0_tx_rst_ack_n_reset_n),                              //  output,    width = 1,                     o_p0_tx_rst_ack_n.reset_n
		.o_p0_ereset_n                      (hssi_ss_1_o_p0_ereset_n_reset),                                    //  output,    width = 1,                         o_p0_ereset_n.reset_n
		.i_clk_ref                          (hssi_ss_1_i_clk_ref_clk),                                          //   input,    width = 2,                             i_clk_ref.clk
		.i_p0_clk_tx_tod                    (hssi_ss_1_o_p0_clk_tx_div_clk),                                    //   input,    width = 1,                       i_p0_clk_tx_tod.clk
		.i_p0_clk_rx_tod                    (hssi_ss_1_o_p0_clk_rec_div_clk_signal),                            //   input,    width = 1,                       i_p0_clk_rx_tod.clk
		.o_p0_clk_pll                       (hssi_ss_1_o_p0_clk_pll_clk),                                       //  output,    width = 1,                          o_p0_clk_pll.clk
		.o_p0_clk_tx_div                    (hssi_ss_1_o_p0_clk_tx_div_clk),                                    //  output,    width = 1,                       o_p0_clk_tx_div.clk
		.o_p0_clk_rec_div64                 (),                                                                 //  output,    width = 1,                    o_p0_clk_rec_div64.clk
		.o_p0_clk_rec_div                   (hssi_ss_1_o_p0_clk_rec_div_clk_signal),                            //  output,    width = 1,                      o_p0_clk_rec_div.clk
		.i_p0_clk_ptp_sample                (sys_manager_ftile_iopll_ptp_sampling_outclk0_clk)                  //   input,    width = 1,                   i_p0_clk_ptp_sample.clk
	);

	ocm ocm (
		.clk        (sys_manager_clk_100_out_clk_clk),     //   input,    width = 1,   clk1.clk
		.address    (mm_interconnect_0_ocm_s1_address),    //   input,   width = 14,     s1.address
		.clken      (mm_interconnect_0_ocm_s1_clken),      //   input,    width = 1,       .clken
		.chipselect (mm_interconnect_0_ocm_s1_chipselect), //   input,    width = 1,       .chipselect
		.write      (mm_interconnect_0_ocm_s1_write),      //   input,    width = 1,       .write
		.readdata   (mm_interconnect_0_ocm_s1_readdata),   //  output,  width = 128,       .readdata
		.writedata  (mm_interconnect_0_ocm_s1_writedata),  //   input,  width = 128,       .writedata
		.byteenable (mm_interconnect_0_ocm_s1_byteenable), //   input,   width = 16,       .byteenable
		.reset      (rst_controller_reset_out_reset),      //   input,    width = 1, reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)   //   input,    width = 1,       .reset_req
	);

	qsfpdd_status_pio qsfpdd_status_pio (
		.clk        (sys_manager_clk_100_out_clk_clk),                   //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_0_qsfpdd_status_pio_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_0_qsfpdd_status_pio_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_0_qsfpdd_status_pio_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_0_qsfpdd_status_pio_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_0_qsfpdd_status_pio_s1_readdata),   //  output,  width = 32,                    .readdata
		.in_port    (qsfpdd_status_pio_external_connection_export),      //   input,   width = 2, external_connection.export
		.irq        (irq_mapper_receiver6_irq)                           //  output,   width = 1,                 irq.irq
	);

	qsfpdd_ctrl_pio_0 sys_ctrl_pio_0 (
		.clk        (sys_manager_clk_100_out_clk_clk),                //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_0_sys_ctrl_pio_0_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_0_sys_ctrl_pio_0_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_0_sys_ctrl_pio_0_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_0_sys_ctrl_pio_0_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_0_sys_ctrl_pio_0_s1_readdata),   //  output,  width = 32,                    .readdata
		.out_port   (qsfpdd_ctrl_pio_0_econ_export)                   //  output,   width = 6, external_connection.export
	);

	clk_ss clk_ss_0 (
		.clk_csr_in_clk_clk                  (clk_csr_in_clk_clk),                    //   input,  width = 1,                  clk_csr_in_clk.clk
		.clk_csr_out_clk_clk                 (clk_ss_0_clk_csr_out_clk_clk),          //  output,  width = 1,                 clk_csr_out_clk.clk
		.clk_dsp_in_clk_clk                  (clk_dsp_in_clk_clk),                    //   input,  width = 1,                  clk_dsp_in_clk.clk
		.clk_dsp_out_clk_clk                 (clk_ss_0_clk_dsp_out_clk_clk),          //  output,  width = 1,                 clk_dsp_out_clk.clk
		.clk_eth_in_clk_clk                  (hssi_ss_1_o_p0_clk_rec_div_clk_signal), //   input,  width = 1,                  clk_eth_in_clk.clk
		.clk_eth_out_clk_clk                 (clk_ss_0_clk_eth_out_clk_clk),          //  output,  width = 1,                 clk_eth_out_clk.clk
		.clk_ftile_402_in_clk_clk            (hssi_ss_1_o_p0_clk_pll_clk),            //   input,  width = 1,            clk_ftile_402_in_clk.clk
		.clk_ftile_402_out_clk_clk           (clk_ss_0_clk_ftile_402_out_clk_clk),    //  output,  width = 1,           clk_ftile_402_out_clk.clk
		.clock_bridge_rec_rx_in_clk_clk      (hssi_ss_1_o_p0_clk_rec_div_clk_signal), //   input,  width = 1,      clock_bridge_rec_rx_in_clk.clk
		.clock_bridge_rec_rx_out_clk_clk     (hssi_ss_1_o_p0_clk_rec_div_clk),        //  output,  width = 1,     clock_bridge_rec_rx_out_clk.clk
		.clock_bridge_rec_rx_out_clk_dup_clk (),                                      //  output,  width = 1, clock_bridge_rec_rx_out_clk_dup.clk
		.ftile_in_clk_clk                    (hssi_ss_1_o_p0_clk_pll_clk),            //   input,  width = 1,                    ftile_in_clk.clk
		.ftile_out_clk_clk                   (ftile_out_clk_clk)                      //  output,  width = 1,                   ftile_out_clk.clk
	);

	ed_synth dfd_subsystem (
		.capture_if_reset_soft_n_rst_soft_n                 (phipps_peak_0_rst_soft_n_dup4_rst_soft_n),                             //   input,    width = 1,        capture_if_reset_soft_n.rst_soft_n
		.capture_if_radio_config_status_radio_config_status (phipps_peak_0_radio_config_status_dup2_radio_config_status),           //   input,   width = 56, capture_if_radio_config_status.radio_config_status
		.lphy_avst_sink_dsp_capture_valid                   (phipps_peak_0_lphy_avst_selctd_cap_intf_valid),                        //   input,    width = 1,     lphy_avst_sink_dsp_capture.valid
		.lphy_avst_sink_dsp_capture_data                    (phipps_peak_0_lphy_avst_selctd_cap_intf_data),                         //   input,   width = 32,                               .data
		.lphy_avst_sink_dsp_capture_channel                 (phipps_peak_0_lphy_avst_selctd_cap_intf_channel),                      //   input,    width = 3,                               .channel
		.dxc_avst_sink_dsp_capture_valid                    (phipps_peak_0_dxc_avst_selctd_cap_intf_valid),                         //   input,    width = 1,      dxc_avst_sink_dsp_capture.valid
		.dxc_avst_sink_dsp_capture_data                     (phipps_peak_0_dxc_avst_selctd_cap_intf_data),                          //   input,   width = 32,                               .data
		.dxc_avst_sink_dsp_capture_channel                  (phipps_peak_0_dxc_avst_selctd_cap_intf_channel),                       //   input,    width = 3,                               .channel
		.interface_sel_data                                 (dfd_subsystem_interface_sel_data),                                     //  output,   width = 32,                  interface_sel.data
		.dsp_in_clk_clk                                     (clk_ss_0_clk_dsp_out_clk_clk),                                         //   input,    width = 1,                     dsp_in_clk.clk
		.eth_in_clk_clk                                     (clk_ss_0_clk_eth_out_clk_clk),                                         //   input,    width = 1,                     eth_in_clk.clk
		.clock_csr_clk                                      (clk_ss_0_clk_csr_out_clk_clk),                                         //   input,    width = 1,                      clock_csr.clk
		.clock_bridge_dspby2_in_clk_clk                     (dfd_subsystem_clock_bridge_dspby2_in_clk_clk),                         //   input,    width = 1,     clock_bridge_dspby2_in_clk.clk
		.ed_synth_h2f_bridge_s0_waitrequest                 (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_waitrequest),   //  output,    width = 1,         ed_synth_h2f_bridge_s0.waitrequest
		.ed_synth_h2f_bridge_s0_readdata                    (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_readdata),      //  output,  width = 512,                               .readdata
		.ed_synth_h2f_bridge_s0_readdatavalid               (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_readdatavalid), //  output,    width = 1,                               .readdatavalid
		.ed_synth_h2f_bridge_s0_burstcount                  (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_burstcount),    //   input,    width = 1,                               .burstcount
		.ed_synth_h2f_bridge_s0_writedata                   (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_writedata),     //   input,  width = 512,                               .writedata
		.ed_synth_h2f_bridge_s0_address                     (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_address),       //   input,   width = 28,                               .address
		.ed_synth_h2f_bridge_s0_write                       (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_write),         //   input,    width = 1,                               .write
		.ed_synth_h2f_bridge_s0_read                        (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_read),          //   input,    width = 1,                               .read
		.ed_synth_h2f_bridge_s0_byteenable                  (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_byteenable),    //   input,   width = 64,                               .byteenable
		.ed_synth_h2f_bridge_s0_debugaccess                 (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_debugaccess),   //   input,    width = 1,                               .debugaccess
		.h2f_lw_bridge_s0_waitrequest                       (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_waitrequest),         //  output,    width = 1,               h2f_lw_bridge_s0.waitrequest
		.h2f_lw_bridge_s0_readdata                          (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_readdata),            //  output,   width = 32,                               .readdata
		.h2f_lw_bridge_s0_readdatavalid                     (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_readdatavalid),       //  output,    width = 1,                               .readdatavalid
		.h2f_lw_bridge_s0_burstcount                        (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_burstcount),          //   input,    width = 1,                               .burstcount
		.h2f_lw_bridge_s0_writedata                         (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_writedata),           //   input,   width = 32,                               .writedata
		.h2f_lw_bridge_s0_address                           (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_address),             //   input,   width = 13,                               .address
		.h2f_lw_bridge_s0_write                             (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_write),               //   input,    width = 1,                               .write
		.h2f_lw_bridge_s0_read                              (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_read),                //   input,    width = 1,                               .read
		.h2f_lw_bridge_s0_byteenable                        (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_byteenable),          //   input,    width = 4,                               .byteenable
		.h2f_lw_bridge_s0_debugaccess                       (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_debugaccess),         //   input,    width = 1,                               .debugaccess
		.dsp_in_reset_reset_n                               (~rst_ss_0_dsp_rst_cntrl_reset_out_reset),                              //   input,    width = 1,                   dsp_in_reset.reset_n
		.eth_in_reset_reset_n                               (~rst_ss_0_eth_rst_cntrl_reset_out_reset),                              //   input,    width = 1,                   eth_in_reset.reset_n
		.reset_csr_reset_n                                  (rst_ss_0_rst_csr_out_reset_reset),                                     //   input,    width = 1,                      reset_csr.reset_n
		.wr_msgdma_0_csr_irq_irq                            ()                                                                      //  output,    width = 1,            wr_msgdma_0_csr_irq.irq
	);

	dma_subsystem dma_subsys (
		.acp_bridge_in_clk_clk                                                        (dma_subsys_acp_bridge_in_clk_clk),                                                        //  output,    width = 1,                                                acp_bridge_in_clk.clk
		.dma_clk_100_in_clk_clk                                                       (sys_manager_clk_100_out_clk_clk),                                                         //   input,    width = 1,                                               dma_clk_100_in_clk.clk
		.dma_clk_out_bridge_0_out_clk_clk                                             (dma_subsys_dma_clk_out_bridge_0_out_clk_clk),                                             //  output,    width = 1,                                     dma_clk_out_bridge_0_out_clk.clk
		.dma_rst_100_in_reset_reset                                                   (rst_controller_reset_out_reset),                                                          //   input,    width = 1,                                             dma_rst_100_in_reset.reset
		.dma_ss_master_m0_waitrequest                                                 (dma_subsys_dma_ss_master_m0_waitrequest),                                                 //   input,    width = 1,                                                 dma_ss_master_m0.waitrequest
		.dma_ss_master_m0_readdata                                                    (dma_subsys_dma_ss_master_m0_readdata),                                                    //   input,  width = 512,                                                                 .readdata
		.dma_ss_master_m0_readdatavalid                                               (dma_subsys_dma_ss_master_m0_readdatavalid),                                               //   input,    width = 1,                                                                 .readdatavalid
		.dma_ss_master_m0_response                                                    (dma_subsys_dma_ss_master_m0_response),                                                    //   input,    width = 2,                                                                 .response
		.dma_ss_master_m0_burstcount                                                  (dma_subsys_dma_ss_master_m0_burstcount),                                                  //  output,    width = 5,                                                                 .burstcount
		.dma_ss_master_m0_writedata                                                   (dma_subsys_dma_ss_master_m0_writedata),                                                   //  output,  width = 512,                                                                 .writedata
		.dma_ss_master_m0_address                                                     (dma_subsys_dma_ss_master_m0_address),                                                     //  output,   width = 37,                                                                 .address
		.dma_ss_master_m0_write                                                       (dma_subsys_dma_ss_master_m0_write),                                                       //  output,    width = 1,                                                                 .write
		.dma_ss_master_m0_read                                                        (dma_subsys_dma_ss_master_m0_read),                                                        //  output,    width = 1,                                                                 .read
		.dma_ss_master_m0_byteenable                                                  (dma_subsys_dma_ss_master_m0_byteenable),                                                  //  output,   width = 64,                                                                 .byteenable
		.dma_ss_master_m0_debugaccess                                                 (dma_subsys_dma_ss_master_m0_debugaccess),                                                 //  output,    width = 1,                                                                 .debugaccess
		.dma_ss_master_m0_writeresponsevalid                                          (dma_subsys_dma_ss_master_m0_writeresponsevalid),                                          //   input,    width = 1,                                                                 .writeresponsevalid
		.ext_hps_m_master_windowed_slave_address                                      (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_address),                    //   input,   width = 30,                                  ext_hps_m_master_windowed_slave.address
		.ext_hps_m_master_windowed_slave_read                                         (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_read),                       //   input,    width = 1,                                                                 .read
		.ext_hps_m_master_windowed_slave_readdata                                     (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_readdata),                   //  output,   width = 32,                                                                 .readdata
		.ext_hps_m_master_windowed_slave_write                                        (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_write),                      //   input,    width = 1,                                                                 .write
		.ext_hps_m_master_windowed_slave_writedata                                    (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_writedata),                  //   input,   width = 32,                                                                 .writedata
		.ext_hps_m_master_windowed_slave_readdatavalid                                (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_readdatavalid),              //  output,    width = 1,                                                                 .readdatavalid
		.ext_hps_m_master_windowed_slave_waitrequest                                  (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_waitrequest),                //  output,    width = 1,                                                                 .waitrequest
		.ext_hps_m_master_windowed_slave_byteenable                                   (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_byteenable),                 //   input,    width = 4,                                                                 .byteenable
		.ext_hps_m_master_windowed_slave_burstcount                                   (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_burstcount),                 //   input,    width = 1,                                                                 .burstcount
		.ext_hps_m_master_expanded_master_address                                     (dma_subsys_ext_hps_m_master_expanded_master_address),                                     //  output,   width = 37,                                 ext_hps_m_master_expanded_master.address
		.ext_hps_m_master_expanded_master_read                                        (dma_subsys_ext_hps_m_master_expanded_master_read),                                        //  output,    width = 1,                                                                 .read
		.ext_hps_m_master_expanded_master_waitrequest                                 (dma_subsys_ext_hps_m_master_expanded_master_waitrequest),                                 //   input,    width = 1,                                                                 .waitrequest
		.ext_hps_m_master_expanded_master_readdata                                    (dma_subsys_ext_hps_m_master_expanded_master_readdata),                                    //   input,   width = 32,                                                                 .readdata
		.ext_hps_m_master_expanded_master_write                                       (dma_subsys_ext_hps_m_master_expanded_master_write),                                       //  output,    width = 1,                                                                 .write
		.ext_hps_m_master_expanded_master_writedata                                   (dma_subsys_ext_hps_m_master_expanded_master_writedata),                                   //  output,   width = 32,                                                                 .writedata
		.ext_hps_m_master_expanded_master_readdatavalid                               (dma_subsys_ext_hps_m_master_expanded_master_readdatavalid),                               //   input,    width = 1,                                                                 .readdatavalid
		.ext_hps_m_master_expanded_master_byteenable                                  (dma_subsys_ext_hps_m_master_expanded_master_byteenable),                                  //  output,    width = 4,                                                                 .byteenable
		.ext_hps_m_master_expanded_master_burstcount                                  (dma_subsys_ext_hps_m_master_expanded_master_burstcount),                                  //  output,    width = 1,                                                                 .burstcount
		.oclk_pll_port8_in_clk_clk                                                    (clk_ss_0_clk_ftile_402_out_clk_clk),                                                      //   input,    width = 1,                                            oclk_pll_port8_in_clk.clk
		.rx_dma_reset_bridge_0_in_reset_reset_n                                       (sys_manager_dma_subsys_port0_rx_dma_resetn_out_reset_reset),                              //   input,    width = 1,                                   rx_dma_reset_bridge_0_in_reset.reset_n
		.rx_dma_reset_bridge_1_in_reset_reset_n                                       (sys_manager_dma_subsys_port1_rx_dma_resetn_out_reset_reset),                              //   input,    width = 1,                                   rx_dma_reset_bridge_1_in_reset.reset_n
		.subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset_reset_n                    (dma_subsys_subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset_reset),                      //  output,    width = 1,                subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset.reset_n
		.ninit_done_reset                                                             (dma_subsys_ninit_done_reset),                                                             //   input,    width = 1,                                                       ninit_done.reset
		.dma_subsys_port8_csr_waitrequest                                             (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_waitrequest),                           //  output,    width = 1,                                             dma_subsys_port8_csr.waitrequest
		.dma_subsys_port8_csr_readdata                                                (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_readdata),                              //  output,   width = 32,                                                                 .readdata
		.dma_subsys_port8_csr_readdatavalid                                           (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_readdatavalid),                         //  output,    width = 1,                                                                 .readdatavalid
		.dma_subsys_port8_csr_burstcount                                              (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_burstcount),                            //   input,    width = 1,                                                                 .burstcount
		.dma_subsys_port8_csr_writedata                                               (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_writedata),                             //   input,   width = 32,                                                                 .writedata
		.dma_subsys_port8_csr_address                                                 (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_address),                               //   input,    width = 8,                                                                 .address
		.dma_subsys_port8_csr_write                                                   (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_write),                                 //   input,    width = 1,                                                                 .write
		.dma_subsys_port8_csr_read                                                    (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_read),                                  //   input,    width = 1,                                                                 .read
		.dma_subsys_port8_csr_byteenable                                              (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_byteenable),                            //   input,    width = 4,                                                                 .byteenable
		.dma_subsys_port8_csr_debugaccess                                             (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_debugaccess),                           //   input,    width = 1,                                                                 .debugaccess
		.dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_startofpacket                  (phipps_peak_0_ecpri_ext_source_startofpacket),                                            //   input,    width = 1,                    dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin.startofpacket
		.dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_valid                          (phipps_peak_0_ecpri_ext_source_valid),                                                    //   input,    width = 1,                                                                 .valid
		.dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_endofpacket                    (phipps_peak_0_ecpri_ext_source_endofpacket),                                              //   input,    width = 1,                                                                 .endofpacket
		.dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_data                           (phipps_peak_0_ecpri_ext_source_data),                                                     //   input,   width = 64,                                                                 .data
		.dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_empty                          (phipps_peak_0_ecpri_ext_source_empty),                                                    //   input,    width = 3,                                                                 .empty
		.dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_error                          (phipps_peak_0_ecpri_ext_source_error),                                                    //   input,    width = 6,                                                                 .error
		.dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_valid            (dma_subsys_dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_valid),            //   input,    width = 1,      dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts.valid
		.dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_data             (dma_subsys_dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_data),             //   input,   width = 96,                                                                 .data
		.dma_subsys_port8_rx_dma_ch1_irq_irq                                          (irq_mapper_receiver2_irq),                                                                //  output,    width = 1,                                  dma_subsys_port8_rx_dma_ch1_irq.irq
		.dma_subsys_port8_ts_chs_compl_0_clk_bus_in_clk                               (clk_ss_0_clk_ftile_402_out_clk_clk),                                                      //   input,    width = 1,                       dma_subsys_port8_ts_chs_compl_0_clk_bus_in.clk
		.dma_subsys_port8_ts_chs_compl_0_rst_bus_in_reset                             (ts_chs_compl_0_rst_bus_in_reset),                                                         //   input,    width = 1,                       dma_subsys_port8_ts_chs_compl_0_rst_bus_in.reset
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_valid            (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_valid),            //   input,    width = 1,      dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts.valid
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_fingerprint      (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_fingerprint),      //   input,   width = 20,                                                                 .fingerprint
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_data             (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_data),             //   input,   width = 96,                                                                 .data
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready           (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready),           //   input,    width = 1,     dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st.ready
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket   (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket),   //  output,    width = 1,                                                                 .startofpacket
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid           (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid),           //  output,    width = 1,                                                                 .valid
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket     (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket),     //  output,    width = 1,                                                                 .endofpacket
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data            (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data),            //  output,   width = 64,                                                                 .data
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty           (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty),           //  output,    width = 3,                                                                 .empty
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error           (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error),           //  output,    width = 1,                                                                 .error
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_valid       (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_valid),       //  output,    width = 1, dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req.valid
		.dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_fingerprint (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_fingerprint), //  output,   width = 20,                                                                 .fingerprint
		.dma_subsys_port8_tx_dma_ch1_irq_irq                                          (irq_mapper_receiver3_irq)                                                                 //  output,    width = 1,                                  dma_subsys_port8_tx_dma_ch1_irq.irq
	);

	hps_sub_sys hps_sub_sys (
		.acp_0_clock_clk                           (dma_subsys_acp_bridge_in_clk_clk),                                   //   input,    width = 1,                  acp_0_clock.clk
		.acp_0_reset_reset                         (rst_controller_001_reset_out_reset),                                 //   input,    width = 1,                  acp_0_reset.reset
		.acp_0_csr_clock_clk                       (sys_manager_clk_100_out_clk_clk),                                    //   input,    width = 1,              acp_0_csr_clock.clk
		.acp_0_csr_reset_reset                     (rst_controller_reset_out_reset),                                     //   input,    width = 1,              acp_0_csr_reset.reset
		.acp_0_csr_address                         (mm_interconnect_1_hps_sub_sys_acp_0_csr_address),                    //   input,    width = 1,                    acp_0_csr.address
		.acp_0_csr_read                            (mm_interconnect_1_hps_sub_sys_acp_0_csr_read),                       //   input,    width = 1,                             .read
		.acp_0_csr_write                           (mm_interconnect_1_hps_sub_sys_acp_0_csr_write),                      //   input,    width = 1,                             .write
		.acp_0_csr_writedata                       (mm_interconnect_1_hps_sub_sys_acp_0_csr_writedata),                  //   input,   width = 32,                             .writedata
		.acp_0_csr_readdata                        (mm_interconnect_1_hps_sub_sys_acp_0_csr_readdata),                   //  output,   width = 32,                             .readdata
		.acp_0_s0_araddr                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_araddr),                      //   input,   width = 37,                     acp_0_s0.araddr
		.acp_0_s0_arburst                          (mm_interconnect_2_hps_sub_sys_acp_0_s0_arburst),                     //   input,    width = 2,                             .arburst
		.acp_0_s0_arcache                          (mm_interconnect_2_hps_sub_sys_acp_0_s0_arcache),                     //   input,    width = 4,                             .arcache
		.acp_0_s0_arid                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_arid),                        //   input,    width = 4,                             .arid
		.acp_0_s0_arlen                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_arlen),                       //   input,    width = 8,                             .arlen
		.acp_0_s0_arlock                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_arlock),                      //   input,    width = 1,                             .arlock
		.acp_0_s0_arprot                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_arprot),                      //   input,    width = 3,                             .arprot
		.acp_0_s0_arready                          (mm_interconnect_2_hps_sub_sys_acp_0_s0_arready),                     //  output,    width = 1,                             .arready
		.acp_0_s0_arsize                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_arsize),                      //   input,    width = 3,                             .arsize
		.acp_0_s0_arvalid                          (mm_interconnect_2_hps_sub_sys_acp_0_s0_arvalid),                     //   input,    width = 1,                             .arvalid
		.acp_0_s0_awaddr                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_awaddr),                      //   input,   width = 37,                             .awaddr
		.acp_0_s0_awburst                          (mm_interconnect_2_hps_sub_sys_acp_0_s0_awburst),                     //   input,    width = 2,                             .awburst
		.acp_0_s0_awcache                          (mm_interconnect_2_hps_sub_sys_acp_0_s0_awcache),                     //   input,    width = 4,                             .awcache
		.acp_0_s0_awid                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_awid),                        //   input,    width = 4,                             .awid
		.acp_0_s0_awlen                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_awlen),                       //   input,    width = 8,                             .awlen
		.acp_0_s0_awlock                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_awlock),                      //   input,    width = 1,                             .awlock
		.acp_0_s0_awprot                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_awprot),                      //   input,    width = 3,                             .awprot
		.acp_0_s0_awready                          (mm_interconnect_2_hps_sub_sys_acp_0_s0_awready),                     //  output,    width = 1,                             .awready
		.acp_0_s0_awsize                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_awsize),                      //   input,    width = 3,                             .awsize
		.acp_0_s0_awvalid                          (mm_interconnect_2_hps_sub_sys_acp_0_s0_awvalid),                     //   input,    width = 1,                             .awvalid
		.acp_0_s0_bid                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_bid),                         //  output,    width = 4,                             .bid
		.acp_0_s0_bready                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_bready),                      //   input,    width = 1,                             .bready
		.acp_0_s0_bresp                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_bresp),                       //  output,    width = 2,                             .bresp
		.acp_0_s0_bvalid                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_bvalid),                      //  output,    width = 1,                             .bvalid
		.acp_0_s0_rdata                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_rdata),                       //  output,  width = 512,                             .rdata
		.acp_0_s0_rid                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_rid),                         //  output,    width = 4,                             .rid
		.acp_0_s0_rlast                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_rlast),                       //  output,    width = 1,                             .rlast
		.acp_0_s0_rready                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_rready),                      //   input,    width = 1,                             .rready
		.acp_0_s0_rresp                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_rresp),                       //  output,    width = 2,                             .rresp
		.acp_0_s0_rvalid                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_rvalid),                      //  output,    width = 1,                             .rvalid
		.acp_0_s0_wdata                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_wdata),                       //   input,  width = 512,                             .wdata
		.acp_0_s0_wlast                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_wlast),                       //   input,    width = 1,                             .wlast
		.acp_0_s0_wready                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_wready),                      //  output,    width = 1,                             .wready
		.acp_0_s0_wstrb                            (mm_interconnect_2_hps_sub_sys_acp_0_s0_wstrb),                       //   input,   width = 64,                             .wstrb
		.acp_0_s0_wvalid                           (mm_interconnect_2_hps_sub_sys_acp_0_s0_wvalid),                      //   input,    width = 1,                             .wvalid
		.agilex_hps_f2h_stm_hw_events_stm_hwevents (agilex_hps_f2h_stm_hw_events_stm_hwevents),                          //   input,   width = 44, agilex_hps_f2h_stm_hw_events.stm_hwevents
		.agilex_hps_h2f_cs_ntrst                   (agilex_hps_h2f_cs_ntrst),                                            //   input,    width = 1,            agilex_hps_h2f_cs.ntrst
		.agilex_hps_h2f_cs_tck                     (agilex_hps_h2f_cs_tck),                                              //   input,    width = 1,                             .tck
		.agilex_hps_h2f_cs_tdi                     (agilex_hps_h2f_cs_tdi),                                              //   input,    width = 1,                             .tdi
		.agilex_hps_h2f_cs_tdo                     (agilex_hps_h2f_cs_tdo),                                              //  output,    width = 1,                             .tdo
		.agilex_hps_h2f_cs_tdoen                   (agilex_hps_h2f_cs_tdoen),                                            //  output,    width = 1,                             .tdoen
		.agilex_hps_h2f_cs_tms                     (agilex_hps_h2f_cs_tms),                                              //   input,    width = 1,                             .tms
		.agilex_hps_hps_io_EMAC1_TX_CLK            (hps_io_EMAC1_TX_CLK),                                                //  output,    width = 1,            agilex_hps_hps_io.EMAC1_TX_CLK
		.agilex_hps_hps_io_EMAC1_TXD0              (hps_io_EMAC1_TXD0),                                                  //  output,    width = 1,                             .EMAC1_TXD0
		.agilex_hps_hps_io_EMAC1_TXD1              (hps_io_EMAC1_TXD1),                                                  //  output,    width = 1,                             .EMAC1_TXD1
		.agilex_hps_hps_io_EMAC1_TXD2              (hps_io_EMAC1_TXD2),                                                  //  output,    width = 1,                             .EMAC1_TXD2
		.agilex_hps_hps_io_EMAC1_TXD3              (hps_io_EMAC1_TXD3),                                                  //  output,    width = 1,                             .EMAC1_TXD3
		.agilex_hps_hps_io_EMAC1_RX_CTL            (hps_io_EMAC1_RX_CTL),                                                //   input,    width = 1,                             .EMAC1_RX_CTL
		.agilex_hps_hps_io_EMAC1_TX_CTL            (hps_io_EMAC1_TX_CTL),                                                //  output,    width = 1,                             .EMAC1_TX_CTL
		.agilex_hps_hps_io_EMAC1_RX_CLK            (hps_io_EMAC1_RX_CLK),                                                //   input,    width = 1,                             .EMAC1_RX_CLK
		.agilex_hps_hps_io_EMAC1_RXD0              (hps_io_EMAC1_RXD0),                                                  //   input,    width = 1,                             .EMAC1_RXD0
		.agilex_hps_hps_io_EMAC1_RXD1              (hps_io_EMAC1_RXD1),                                                  //   input,    width = 1,                             .EMAC1_RXD1
		.agilex_hps_hps_io_EMAC1_RXD2              (hps_io_EMAC1_RXD2),                                                  //   input,    width = 1,                             .EMAC1_RXD2
		.agilex_hps_hps_io_EMAC1_RXD3              (hps_io_EMAC1_RXD3),                                                  //   input,    width = 1,                             .EMAC1_RXD3
		.agilex_hps_hps_io_EMAC1_MDIO              (hps_io_EMAC1_MDIO),                                                  //   inout,    width = 1,                             .EMAC1_MDIO
		.agilex_hps_hps_io_EMAC1_MDC               (hps_io_EMAC1_MDC),                                                   //  output,    width = 1,                             .EMAC1_MDC
		.agilex_hps_hps_io_SDMMC_CMD               (hps_io_SDMMC_CMD),                                                   //   inout,    width = 1,                             .SDMMC_CMD
		.agilex_hps_hps_io_SDMMC_D0                (hps_io_SDMMC_D0),                                                    //   inout,    width = 1,                             .SDMMC_D0
		.agilex_hps_hps_io_SDMMC_D1                (hps_io_SDMMC_D1),                                                    //   inout,    width = 1,                             .SDMMC_D1
		.agilex_hps_hps_io_SDMMC_D2                (hps_io_SDMMC_D2),                                                    //   inout,    width = 1,                             .SDMMC_D2
		.agilex_hps_hps_io_SDMMC_D3                (hps_io_SDMMC_D3),                                                    //   inout,    width = 1,                             .SDMMC_D3
		.agilex_hps_hps_io_SDMMC_D4                (hps_io_SDMMC_D4),                                                    //   inout,    width = 1,                             .SDMMC_D4
		.agilex_hps_hps_io_SDMMC_D5                (hps_io_SDMMC_D5),                                                    //   inout,    width = 1,                             .SDMMC_D5
		.agilex_hps_hps_io_SDMMC_D6                (hps_io_SDMMC_D6),                                                    //   inout,    width = 1,                             .SDMMC_D6
		.agilex_hps_hps_io_SDMMC_D7                (hps_io_SDMMC_D7),                                                    //   inout,    width = 1,                             .SDMMC_D7
		.agilex_hps_hps_io_SDMMC_CCLK              (hps_io_SDMMC_CCLK),                                                  //  output,    width = 1,                             .SDMMC_CCLK
		.agilex_hps_hps_io_SPIM0_CLK               (hps_io_SPIM0_CLK),                                                   //  output,    width = 1,                             .SPIM0_CLK
		.agilex_hps_hps_io_SPIM0_MOSI              (hps_io_SPIM0_MOSI),                                                  //  output,    width = 1,                             .SPIM0_MOSI
		.agilex_hps_hps_io_SPIM0_MISO              (hps_io_SPIM0_MISO),                                                  //   input,    width = 1,                             .SPIM0_MISO
		.agilex_hps_hps_io_SPIM0_SS0_N             (hps_io_SPIM0_SS0_N),                                                 //  output,    width = 1,                             .SPIM0_SS0_N
		.agilex_hps_hps_io_SPIM1_CLK               (hps_io_SPIM1_CLK),                                                   //  output,    width = 1,                             .SPIM1_CLK
		.agilex_hps_hps_io_SPIM1_MOSI              (hps_io_SPIM1_MOSI),                                                  //  output,    width = 1,                             .SPIM1_MOSI
		.agilex_hps_hps_io_SPIM1_MISO              (hps_io_SPIM1_MISO),                                                  //   input,    width = 1,                             .SPIM1_MISO
		.agilex_hps_hps_io_SPIM1_SS0_N             (hps_io_SPIM1_SS0_N),                                                 //  output,    width = 1,                             .SPIM1_SS0_N
		.agilex_hps_hps_io_SPIM1_SS1_N             (hps_io_SPIM1_SS1_N),                                                 //  output,    width = 1,                             .SPIM1_SS1_N
		.agilex_hps_hps_io_UART1_RX                (hps_io_UART1_RX),                                                    //   input,    width = 1,                             .UART1_RX
		.agilex_hps_hps_io_UART1_TX                (hps_io_UART1_TX),                                                    //  output,    width = 1,                             .UART1_TX
		.agilex_hps_hps_io_I2C1_SDA                (hps_io_I2C1_SDA),                                                    //   inout,    width = 1,                             .I2C1_SDA
		.agilex_hps_hps_io_I2C1_SCL                (hps_io_I2C1_SCL),                                                    //   inout,    width = 1,                             .I2C1_SCL
		.agilex_hps_hps_io_hps_osc_clk             (hps_io_hps_osc_clk),                                                 //   input,    width = 1,                             .hps_osc_clk
		.agilex_hps_hps_io_gpio0_io11              (hps_io_gpio0_io11),                                                  //   inout,    width = 1,                             .gpio0_io11
		.agilex_hps_hps_io_gpio0_io12              (hps_io_gpio0_io12),                                                  //   inout,    width = 1,                             .gpio0_io12
		.agilex_hps_hps_io_gpio0_io13              (hps_io_gpio0_io13),                                                  //   inout,    width = 1,                             .gpio0_io13
		.agilex_hps_hps_io_gpio0_io14              (hps_io_gpio0_io14),                                                  //   inout,    width = 1,                             .gpio0_io14
		.agilex_hps_hps_io_gpio0_io15              (hps_io_gpio0_io15),                                                  //   inout,    width = 1,                             .gpio0_io15
		.agilex_hps_hps_io_gpio0_io16              (hps_io_gpio0_io16),                                                  //   inout,    width = 1,                             .gpio0_io16
		.agilex_hps_hps_io_gpio0_io17              (hps_io_gpio0_io17),                                                  //   inout,    width = 1,                             .gpio0_io17
		.agilex_hps_hps_io_gpio0_io18              (hps_io_gpio0_io18),                                                  //   inout,    width = 1,                             .gpio0_io18
		.agilex_hps_hps_io_gpio1_io16              (hps_io_gpio1_io16),                                                  //   inout,    width = 1,                             .gpio1_io16
		.agilex_hps_hps_io_gpio1_io17              (hps_io_gpio1_io17),                                                  //   inout,    width = 1,                             .gpio1_io17
		.agilex_hps_h2f_reset_reset                (agilex_hps_h2f_reset_reset),                                         //  output,    width = 1,         agilex_hps_h2f_reset.reset
		.agilex_hps_h2f_axi_clock_clk              (sys_manager_clk_100_out_clk_clk),                                    //   input,    width = 1,     agilex_hps_h2f_axi_clock.clk
		.agilex_hps_h2f_axi_reset_reset_n          (~rst_controller_reset_out_reset),                                    //   input,    width = 1,     agilex_hps_h2f_axi_reset.reset_n
		.agilex_hps_h2f_axi_master_awid            (hps_sub_sys_agilex_hps_h2f_axi_master_awid),                         //  output,    width = 4,    agilex_hps_h2f_axi_master.awid
		.agilex_hps_h2f_axi_master_awaddr          (hps_sub_sys_agilex_hps_h2f_axi_master_awaddr),                       //  output,   width = 32,                             .awaddr
		.agilex_hps_h2f_axi_master_awlen           (hps_sub_sys_agilex_hps_h2f_axi_master_awlen),                        //  output,    width = 8,                             .awlen
		.agilex_hps_h2f_axi_master_awsize          (hps_sub_sys_agilex_hps_h2f_axi_master_awsize),                       //  output,    width = 3,                             .awsize
		.agilex_hps_h2f_axi_master_awburst         (hps_sub_sys_agilex_hps_h2f_axi_master_awburst),                      //  output,    width = 2,                             .awburst
		.agilex_hps_h2f_axi_master_awlock          (hps_sub_sys_agilex_hps_h2f_axi_master_awlock),                       //  output,    width = 1,                             .awlock
		.agilex_hps_h2f_axi_master_awcache         (hps_sub_sys_agilex_hps_h2f_axi_master_awcache),                      //  output,    width = 4,                             .awcache
		.agilex_hps_h2f_axi_master_awprot          (hps_sub_sys_agilex_hps_h2f_axi_master_awprot),                       //  output,    width = 3,                             .awprot
		.agilex_hps_h2f_axi_master_awvalid         (hps_sub_sys_agilex_hps_h2f_axi_master_awvalid),                      //  output,    width = 1,                             .awvalid
		.agilex_hps_h2f_axi_master_awready         (hps_sub_sys_agilex_hps_h2f_axi_master_awready),                      //   input,    width = 1,                             .awready
		.agilex_hps_h2f_axi_master_wdata           (hps_sub_sys_agilex_hps_h2f_axi_master_wdata),                        //  output,  width = 128,                             .wdata
		.agilex_hps_h2f_axi_master_wstrb           (hps_sub_sys_agilex_hps_h2f_axi_master_wstrb),                        //  output,   width = 16,                             .wstrb
		.agilex_hps_h2f_axi_master_wlast           (hps_sub_sys_agilex_hps_h2f_axi_master_wlast),                        //  output,    width = 1,                             .wlast
		.agilex_hps_h2f_axi_master_wvalid          (hps_sub_sys_agilex_hps_h2f_axi_master_wvalid),                       //  output,    width = 1,                             .wvalid
		.agilex_hps_h2f_axi_master_wready          (hps_sub_sys_agilex_hps_h2f_axi_master_wready),                       //   input,    width = 1,                             .wready
		.agilex_hps_h2f_axi_master_bid             (hps_sub_sys_agilex_hps_h2f_axi_master_bid),                          //   input,    width = 4,                             .bid
		.agilex_hps_h2f_axi_master_bresp           (hps_sub_sys_agilex_hps_h2f_axi_master_bresp),                        //   input,    width = 2,                             .bresp
		.agilex_hps_h2f_axi_master_bvalid          (hps_sub_sys_agilex_hps_h2f_axi_master_bvalid),                       //   input,    width = 1,                             .bvalid
		.agilex_hps_h2f_axi_master_bready          (hps_sub_sys_agilex_hps_h2f_axi_master_bready),                       //  output,    width = 1,                             .bready
		.agilex_hps_h2f_axi_master_arid            (hps_sub_sys_agilex_hps_h2f_axi_master_arid),                         //  output,    width = 4,                             .arid
		.agilex_hps_h2f_axi_master_araddr          (hps_sub_sys_agilex_hps_h2f_axi_master_araddr),                       //  output,   width = 32,                             .araddr
		.agilex_hps_h2f_axi_master_arlen           (hps_sub_sys_agilex_hps_h2f_axi_master_arlen),                        //  output,    width = 8,                             .arlen
		.agilex_hps_h2f_axi_master_arsize          (hps_sub_sys_agilex_hps_h2f_axi_master_arsize),                       //  output,    width = 3,                             .arsize
		.agilex_hps_h2f_axi_master_arburst         (hps_sub_sys_agilex_hps_h2f_axi_master_arburst),                      //  output,    width = 2,                             .arburst
		.agilex_hps_h2f_axi_master_arlock          (hps_sub_sys_agilex_hps_h2f_axi_master_arlock),                       //  output,    width = 1,                             .arlock
		.agilex_hps_h2f_axi_master_arcache         (hps_sub_sys_agilex_hps_h2f_axi_master_arcache),                      //  output,    width = 4,                             .arcache
		.agilex_hps_h2f_axi_master_arprot          (hps_sub_sys_agilex_hps_h2f_axi_master_arprot),                       //  output,    width = 3,                             .arprot
		.agilex_hps_h2f_axi_master_arvalid         (hps_sub_sys_agilex_hps_h2f_axi_master_arvalid),                      //  output,    width = 1,                             .arvalid
		.agilex_hps_h2f_axi_master_arready         (hps_sub_sys_agilex_hps_h2f_axi_master_arready),                      //   input,    width = 1,                             .arready
		.agilex_hps_h2f_axi_master_rid             (hps_sub_sys_agilex_hps_h2f_axi_master_rid),                          //   input,    width = 4,                             .rid
		.agilex_hps_h2f_axi_master_rdata           (hps_sub_sys_agilex_hps_h2f_axi_master_rdata),                        //   input,  width = 128,                             .rdata
		.agilex_hps_h2f_axi_master_rresp           (hps_sub_sys_agilex_hps_h2f_axi_master_rresp),                        //   input,    width = 2,                             .rresp
		.agilex_hps_h2f_axi_master_rlast           (hps_sub_sys_agilex_hps_h2f_axi_master_rlast),                        //   input,    width = 1,                             .rlast
		.agilex_hps_h2f_axi_master_rvalid          (hps_sub_sys_agilex_hps_h2f_axi_master_rvalid),                       //   input,    width = 1,                             .rvalid
		.agilex_hps_h2f_axi_master_rready          (hps_sub_sys_agilex_hps_h2f_axi_master_rready),                       //  output,    width = 1,                             .rready
		.agilex_hps_h2f_lw_axi_clock_clk           (sys_manager_clk_100_out_clk_clk),                                    //   input,    width = 1,  agilex_hps_h2f_lw_axi_clock.clk
		.agilex_hps_h2f_lw_axi_reset_reset_n       (~rst_controller_reset_out_reset),                                    //   input,    width = 1,  agilex_hps_h2f_lw_axi_reset.reset_n
		.agilex_hps_h2f_lw_axi_master_awid         (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awid),                      //  output,    width = 4, agilex_hps_h2f_lw_axi_master.awid
		.agilex_hps_h2f_lw_axi_master_awaddr       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awaddr),                    //  output,   width = 21,                             .awaddr
		.agilex_hps_h2f_lw_axi_master_awlen        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlen),                     //  output,    width = 8,                             .awlen
		.agilex_hps_h2f_lw_axi_master_awsize       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awsize),                    //  output,    width = 3,                             .awsize
		.agilex_hps_h2f_lw_axi_master_awburst      (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awburst),                   //  output,    width = 2,                             .awburst
		.agilex_hps_h2f_lw_axi_master_awlock       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlock),                    //  output,    width = 1,                             .awlock
		.agilex_hps_h2f_lw_axi_master_awcache      (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awcache),                   //  output,    width = 4,                             .awcache
		.agilex_hps_h2f_lw_axi_master_awprot       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awprot),                    //  output,    width = 3,                             .awprot
		.agilex_hps_h2f_lw_axi_master_awvalid      (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awvalid),                   //  output,    width = 1,                             .awvalid
		.agilex_hps_h2f_lw_axi_master_awready      (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awready),                   //   input,    width = 1,                             .awready
		.agilex_hps_h2f_lw_axi_master_wdata        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wdata),                     //  output,   width = 32,                             .wdata
		.agilex_hps_h2f_lw_axi_master_wstrb        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wstrb),                     //  output,    width = 4,                             .wstrb
		.agilex_hps_h2f_lw_axi_master_wlast        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wlast),                     //  output,    width = 1,                             .wlast
		.agilex_hps_h2f_lw_axi_master_wvalid       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wvalid),                    //  output,    width = 1,                             .wvalid
		.agilex_hps_h2f_lw_axi_master_wready       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wready),                    //   input,    width = 1,                             .wready
		.agilex_hps_h2f_lw_axi_master_bid          (hps_sub_sys_agilex_hps_h2f_lw_axi_master_bid),                       //   input,    width = 4,                             .bid
		.agilex_hps_h2f_lw_axi_master_bresp        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_bresp),                     //   input,    width = 2,                             .bresp
		.agilex_hps_h2f_lw_axi_master_bvalid       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_bvalid),                    //   input,    width = 1,                             .bvalid
		.agilex_hps_h2f_lw_axi_master_bready       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_bready),                    //  output,    width = 1,                             .bready
		.agilex_hps_h2f_lw_axi_master_arid         (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arid),                      //  output,    width = 4,                             .arid
		.agilex_hps_h2f_lw_axi_master_araddr       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_araddr),                    //  output,   width = 21,                             .araddr
		.agilex_hps_h2f_lw_axi_master_arlen        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlen),                     //  output,    width = 8,                             .arlen
		.agilex_hps_h2f_lw_axi_master_arsize       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arsize),                    //  output,    width = 3,                             .arsize
		.agilex_hps_h2f_lw_axi_master_arburst      (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arburst),                   //  output,    width = 2,                             .arburst
		.agilex_hps_h2f_lw_axi_master_arlock       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlock),                    //  output,    width = 1,                             .arlock
		.agilex_hps_h2f_lw_axi_master_arcache      (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arcache),                   //  output,    width = 4,                             .arcache
		.agilex_hps_h2f_lw_axi_master_arprot       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arprot),                    //  output,    width = 3,                             .arprot
		.agilex_hps_h2f_lw_axi_master_arvalid      (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arvalid),                   //  output,    width = 1,                             .arvalid
		.agilex_hps_h2f_lw_axi_master_arready      (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arready),                   //   input,    width = 1,                             .arready
		.agilex_hps_h2f_lw_axi_master_rid          (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rid),                       //   input,    width = 4,                             .rid
		.agilex_hps_h2f_lw_axi_master_rdata        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rdata),                     //   input,   width = 32,                             .rdata
		.agilex_hps_h2f_lw_axi_master_rresp        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rresp),                     //   input,    width = 2,                             .rresp
		.agilex_hps_h2f_lw_axi_master_rlast        (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rlast),                     //   input,    width = 1,                             .rlast
		.agilex_hps_h2f_lw_axi_master_rvalid       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rvalid),                    //   input,    width = 1,                             .rvalid
		.agilex_hps_h2f_lw_axi_master_rready       (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rready),                    //  output,    width = 1,                             .rready
		.agilex_hps_f2h_axi_clock_clk              (dma_subsys_dma_clk_out_bridge_0_out_clk_clk),                        //   input,    width = 1,     agilex_hps_f2h_axi_clock.clk
		.agilex_hps_f2h_axi_reset_reset_n          (dma_subsys_subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset_reset), //   input,    width = 1,     agilex_hps_f2h_axi_reset.reset_n
		.agilex_hps_f2h_irq0_irq                   (hps_sub_sys_agilex_hps_f2h_irq0_irq),                                //   input,   width = 32,          agilex_hps_f2h_irq0.irq
		.agilex_hps_f2h_irq1_irq                   (f2h_irq1_irq),                                                       //   input,   width = 32,          agilex_hps_f2h_irq1.irq
		.emif_hps_pll_ref_clk_clk                  (emif_hps_pll_ref_clk_clk),                                           //   input,    width = 1,         emif_hps_pll_ref_clk.clk
		.emif_hps_oct_oct_rzqin                    (emif_hps_oct_oct_rzqin),                                             //   input,    width = 1,                 emif_hps_oct.oct_rzqin
		.emif_hps_mem_mem_ck                       (emif_hps_mem_mem_ck),                                                //  output,    width = 1,                 emif_hps_mem.mem_ck
		.emif_hps_mem_mem_ck_n                     (emif_hps_mem_mem_ck_n),                                              //  output,    width = 1,                             .mem_ck_n
		.emif_hps_mem_mem_a                        (emif_hps_mem_mem_a),                                                 //  output,   width = 17,                             .mem_a
		.emif_hps_mem_mem_act_n                    (emif_hps_mem_mem_act_n),                                             //  output,    width = 1,                             .mem_act_n
		.emif_hps_mem_mem_ba                       (emif_hps_mem_mem_ba),                                                //  output,    width = 2,                             .mem_ba
		.emif_hps_mem_mem_bg                       (emif_hps_mem_mem_bg),                                                //  output,    width = 1,                             .mem_bg
		.emif_hps_mem_mem_cke                      (emif_hps_mem_mem_cke),                                               //  output,    width = 1,                             .mem_cke
		.emif_hps_mem_mem_cs_n                     (emif_hps_mem_mem_cs_n),                                              //  output,    width = 2,                             .mem_cs_n
		.emif_hps_mem_mem_odt                      (emif_hps_mem_mem_odt),                                               //  output,    width = 1,                             .mem_odt
		.emif_hps_mem_mem_reset_n                  (emif_hps_mem_mem_reset_n),                                           //  output,    width = 1,                             .mem_reset_n
		.emif_hps_mem_mem_par                      (emif_hps_mem_mem_par),                                               //  output,    width = 1,                             .mem_par
		.emif_hps_mem_mem_alert_n                  (emif_hps_mem_mem_alert_n),                                           //   input,    width = 1,                             .mem_alert_n
		.emif_hps_mem_mem_dqs                      (emif_hps_mem_mem_dqs),                                               //   inout,    width = 9,                             .mem_dqs
		.emif_hps_mem_mem_dqs_n                    (emif_hps_mem_mem_dqs_n),                                             //   inout,    width = 9,                             .mem_dqs_n
		.emif_hps_mem_mem_dq                       (emif_hps_mem_mem_dq),                                                //   inout,   width = 72,                             .mem_dq
		.emif_hps_mem_mem_dbi_n                    (emif_hps_mem_mem_dbi_n)                                              //   inout,    width = 9,                             .mem_dbi_n
	);

	j204c_f_rx_tx_ip j204c_f_rx_tx_ip (
		.intel_jesd204c_f_reconfig_xcvr_address        (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_address),     //   input,   width = 21,         intel_jesd204c_f_reconfig_xcvr.address
		.intel_jesd204c_f_reconfig_xcvr_read           (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_read),        //   input,    width = 1,                                       .read
		.intel_jesd204c_f_reconfig_xcvr_write          (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_write),       //   input,    width = 1,                                       .write
		.intel_jesd204c_f_reconfig_xcvr_writedata      (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_writedata),   //   input,   width = 32,                                       .writedata
		.intel_jesd204c_f_reconfig_xcvr_readdata       (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_readdata),    //  output,   width = 32,                                       .readdata
		.intel_jesd204c_f_reconfig_xcvr_waitrequest    (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_waitrequest), //  output,    width = 1,                                       .waitrequest
		.intel_jesd204c_f_reconfig_xcvr_byteenable     (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_byteenable),  //   input,    width = 4,                                       .byteenable
		.intel_jesd204c_f_j204c_tx_rst_ack_n_export    (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_rst_ack_n_export),                   //  output,    width = 1,    intel_jesd204c_f_j204c_tx_rst_ack_n.export
		.intel_jesd204c_f_j204c_txlclk_ctrl_export     (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_txlclk_ctrl_export),                    //   input,    width = 1,     intel_jesd204c_f_j204c_txlclk_ctrl.export
		.intel_jesd204c_f_j204c_txfclk_ctrl_export     (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_txfclk_ctrl_export),                    //   input,    width = 1,     intel_jesd204c_f_j204c_txfclk_ctrl.export
		.intel_jesd204c_f_j204c_tx_avs_chipselect      (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_chipselect),   //   input,    width = 1,          intel_jesd204c_f_j204c_tx_avs.chipselect
		.intel_jesd204c_f_j204c_tx_avs_address         (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_address),      //   input,   width = 10,                                       .address
		.intel_jesd204c_f_j204c_tx_avs_read            (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_read),         //   input,    width = 1,                                       .read
		.intel_jesd204c_f_j204c_tx_avs_readdata        (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_readdata),     //  output,   width = 32,                                       .readdata
		.intel_jesd204c_f_j204c_tx_avs_waitrequest     (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_waitrequest),  //  output,    width = 1,                                       .waitrequest
		.intel_jesd204c_f_j204c_tx_avs_write           (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_write),        //   input,    width = 1,                                       .write
		.intel_jesd204c_f_j204c_tx_avs_writedata       (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_writedata),    //   input,   width = 32,                                       .writedata
		.intel_jesd204c_f_j204c_tx_avst_data           (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avst_data),                          //   input,  width = 512,         intel_jesd204c_f_j204c_tx_avst.data
		.intel_jesd204c_f_j204c_tx_avst_valid          (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avst_valid),                         //   input,    width = 1,                                       .valid
		.intel_jesd204c_f_j204c_tx_avst_ready          (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avst_ready),                         //  output,    width = 1,                                       .ready
		.intel_jesd204c_f_j204c_tx_avst_control_export (),                                                                              //   input,    width = 1, intel_jesd204c_f_j204c_tx_avst_control.export
		.intel_jesd204c_f_j204c_tx_cmd_data            (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_cmd_data),                           //   input,   width = 48,          intel_jesd204c_f_j204c_tx_cmd.data
		.intel_jesd204c_f_j204c_tx_cmd_valid           (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_cmd_valid),                          //   input,    width = 1,                                       .valid
		.intel_jesd204c_f_j204c_tx_cmd_ready           (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_cmd_ready),                          //  output,    width = 1,                                       .ready
		.intel_jesd204c_f_j204c_tx_sysref_export       (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_sysref_export),                      //   input,    width = 1,       intel_jesd204c_f_j204c_tx_sysref.export
		.intel_jesd204c_f_j204c_tx_csr_l_export        (),                                                                              //  output,    width = 4,        intel_jesd204c_f_j204c_tx_csr_l.export
		.intel_jesd204c_f_j204c_tx_csr_f_export        (),                                                                              //  output,    width = 8,        intel_jesd204c_f_j204c_tx_csr_f.export
		.intel_jesd204c_f_j204c_tx_csr_m_export        (),                                                                              //  output,    width = 8,        intel_jesd204c_f_j204c_tx_csr_m.export
		.intel_jesd204c_f_j204c_tx_csr_cs_export       (),                                                                              //  output,    width = 2,       intel_jesd204c_f_j204c_tx_csr_cs.export
		.intel_jesd204c_f_j204c_tx_csr_n_export        (),                                                                              //  output,    width = 5,        intel_jesd204c_f_j204c_tx_csr_n.export
		.intel_jesd204c_f_j204c_tx_csr_np_export       (),                                                                              //  output,    width = 5,       intel_jesd204c_f_j204c_tx_csr_np.export
		.intel_jesd204c_f_j204c_tx_csr_s_export        (),                                                                              //  output,    width = 5,        intel_jesd204c_f_j204c_tx_csr_s.export
		.intel_jesd204c_f_j204c_tx_csr_hd_export       (),                                                                              //  output,    width = 1,       intel_jesd204c_f_j204c_tx_csr_hd.export
		.intel_jesd204c_f_j204c_tx_csr_cf_export       (),                                                                              //  output,    width = 5,       intel_jesd204c_f_j204c_tx_csr_cf.export
		.intel_jesd204c_f_j204c_tx_csr_e_export        (),                                                                              //  output,    width = 8,        intel_jesd204c_f_j204c_tx_csr_e.export
		.intel_jesd204c_f_j204c_tx_int_irq             (),                                                                              //  output,    width = 1,          intel_jesd204c_f_j204c_tx_int.irq
		.intel_jesd204c_f_j204c_rx_avs_chipselect      (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_chipselect),   //   input,    width = 1,          intel_jesd204c_f_j204c_rx_avs.chipselect
		.intel_jesd204c_f_j204c_rx_avs_address         (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_address),      //   input,   width = 10,                                       .address
		.intel_jesd204c_f_j204c_rx_avs_read            (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_read),         //   input,    width = 1,                                       .read
		.intel_jesd204c_f_j204c_rx_avs_readdata        (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_readdata),     //  output,   width = 32,                                       .readdata
		.intel_jesd204c_f_j204c_rx_avs_waitrequest     (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_waitrequest),  //  output,    width = 1,                                       .waitrequest
		.intel_jesd204c_f_j204c_rx_avs_write           (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_write),        //   input,    width = 1,                                       .write
		.intel_jesd204c_f_j204c_rx_avs_writedata       (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_writedata),    //   input,   width = 32,                                       .writedata
		.intel_jesd204c_f_j204c_rx_int_irq             (),                                                                              //  output,    width = 1,          intel_jesd204c_f_j204c_rx_int.irq
		.intel_jesd204c_f_j204c_rx_csr_l_export        (),                                                                              //  output,    width = 4,        intel_jesd204c_f_j204c_rx_csr_l.export
		.intel_jesd204c_f_j204c_rx_csr_f_export        (),                                                                              //  output,    width = 8,        intel_jesd204c_f_j204c_rx_csr_f.export
		.intel_jesd204c_f_j204c_rx_csr_m_export        (),                                                                              //  output,    width = 8,        intel_jesd204c_f_j204c_rx_csr_m.export
		.intel_jesd204c_f_j204c_rx_csr_cs_export       (),                                                                              //  output,    width = 2,       intel_jesd204c_f_j204c_rx_csr_cs.export
		.intel_jesd204c_f_j204c_rx_csr_n_export        (),                                                                              //  output,    width = 5,        intel_jesd204c_f_j204c_rx_csr_n.export
		.intel_jesd204c_f_j204c_rx_csr_np_export       (),                                                                              //  output,    width = 5,       intel_jesd204c_f_j204c_rx_csr_np.export
		.intel_jesd204c_f_j204c_rx_csr_s_export        (),                                                                              //  output,    width = 5,        intel_jesd204c_f_j204c_rx_csr_s.export
		.intel_jesd204c_f_j204c_rx_csr_hd_export       (),                                                                              //  output,    width = 1,       intel_jesd204c_f_j204c_rx_csr_hd.export
		.intel_jesd204c_f_j204c_rx_csr_cf_export       (),                                                                              //  output,    width = 5,       intel_jesd204c_f_j204c_rx_csr_cf.export
		.intel_jesd204c_f_j204c_rx_csr_e_export        (),                                                                              //  output,    width = 8,        intel_jesd204c_f_j204c_rx_csr_e.export
		.intel_jesd204c_f_j204c_rx_csr_testmode_export (),                                                                              //  output,    width = 2, intel_jesd204c_f_j204c_rx_csr_testmode.export
		.intel_jesd204c_f_j204c_rxlclk_ctrl_export     (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rxlclk_ctrl_export),                    //   input,    width = 1,     intel_jesd204c_f_j204c_rxlclk_ctrl.export
		.intel_jesd204c_f_j204c_rxfclk_ctrl_export     (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rxfclk_ctrl_export),                    //   input,    width = 1,     intel_jesd204c_f_j204c_rxfclk_ctrl.export
		.intel_jesd204c_f_j204c_rx_sysref_export       (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_sysref_export),                      //   input,    width = 1,       intel_jesd204c_f_j204c_rx_sysref.export
		.intel_jesd204c_f_j204c_rx_rst_ack_n_export    (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_rst_ack_n_export),                   //  output,    width = 1,    intel_jesd204c_f_j204c_rx_rst_ack_n.export
		.intel_jesd204c_f_j204c_rx_avst_data           (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avst_data),                          //  output,  width = 512,         intel_jesd204c_f_j204c_rx_avst.data
		.intel_jesd204c_f_j204c_rx_avst_valid          (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avst_valid),                         //  output,    width = 1,                                       .valid
		.intel_jesd204c_f_j204c_rx_avst_ready          (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avst_ready),                         //   input,    width = 1,                                       .ready
		.intel_jesd204c_f_j204c_rx_avst_control_export (),                                                                              //  output,    width = 1, intel_jesd204c_f_j204c_rx_avst_control.export
		.intel_jesd204c_f_j204c_rx_cmd_data            (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_cmd_data),                           //  output,   width = 48,          intel_jesd204c_f_j204c_rx_cmd.data
		.intel_jesd204c_f_j204c_rx_cmd_valid           (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_cmd_valid),                          //  output,    width = 1,                                       .valid
		.intel_jesd204c_f_j204c_rx_cmd_ready           (j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_cmd_ready),                          //   input,    width = 1,                                       .ready
		.intel_jesd204c_f_j204c_rx_cmd_par_err_export  (),                                                                              //  output,    width = 8,  intel_jesd204c_f_j204c_rx_cmd_par_err.export
		.intel_jesd204c_f_j204c_rx_sh_lock_export      (),                                                                              //  output,    width = 1,      intel_jesd204c_f_j204c_rx_sh_lock.export
		.intel_jesd204c_f_j204c_rx_emb_lock_export     (),                                                                              //  output,    width = 1,     intel_jesd204c_f_j204c_rx_emb_lock.export
		.intel_jesd204c_f_j204c_rx_crc_err_export      (),                                                                              //  output,    width = 8,      intel_jesd204c_f_j204c_rx_crc_err.export
		.intel_jesd204c_f_tx_serial_data_export        (j204c_f_rx_tx_ip_intel_jesd204c_f_tx_serial_data_export),                       //  output,    width = 8,        intel_jesd204c_f_tx_serial_data.export
		.intel_jesd204c_f_tx_serial_data_n_export      (j204c_f_rx_tx_ip_intel_jesd204c_f_tx_serial_data_n_export),                     //  output,    width = 8,      intel_jesd204c_f_tx_serial_data_n.export
		.intel_jesd204c_f_rx_serial_data_export        (j204c_f_rx_tx_ip_intel_jesd204c_f_rx_serial_data_export),                       //   input,    width = 8,        intel_jesd204c_f_rx_serial_data.export
		.intel_jesd204c_f_rx_serial_data_n_export      (j204c_f_rx_tx_ip_intel_jesd204c_f_rx_serial_data_n_export),                     //   input,    width = 8,      intel_jesd204c_f_rx_serial_data_n.export
		.jesd_link_clk_in_clk_clk                      (j204c_f_rx_tx_ip_jesd_link_clk_in_clk_clk),                                     //   input,    width = 1,                   jesd_link_clk_in_clk.clk
		.mgmt_clk_in_clk_clk                           (sys_manager_clk_100_out_clk_clk),                                               //   input,    width = 1,                        mgmt_clk_in_clk.clk
		.mgmt_reset_in_reset_reset_n                   (~rst_controller_reset_out_reset),                                               //   input,    width = 1,                    mgmt_reset_in_reset.reset_n
		.reset_out1_reset                              (j204c_f_rx_tx_ip_reset_out1_reset),                                             //  output,    width = 1,                             reset_out1.reset
		.reset_out2_reset                              (j204c_f_rx_tx_ip_reset_out2_reset),                                             //  output,    width = 1,                             reset_out2.reset
		.reset_out4_reset                              (j204c_f_rx_tx_ip_reset_out4_reset),                                             //  output,    width = 1,                             reset_out4.reset
		.reset1_dsrt_qual_reset1_dsrt_qual             (j204c_f_rx_tx_ip_reset1_dsrt_qual_reset1_dsrt_qual),                            //   input,    width = 1,                       reset1_dsrt_qual.reset1_dsrt_qual
		.reset2_dsrt_qual_reset2_dsrt_qual             (j204c_f_rx_tx_ip_reset2_dsrt_qual_reset2_dsrt_qual),                            //   input,    width = 1,                       reset2_dsrt_qual.reset2_dsrt_qual
		.reset4_dsrt_qual_reset4_dsrt_qual             (j204c_f_rx_tx_ip_reset4_dsrt_qual_reset4_dsrt_qual),                            //   input,    width = 1,                       reset4_dsrt_qual.reset4_dsrt_qual
		.reset_sequencer_0_av_csr_address              (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_address),           //   input,    width = 8,               reset_sequencer_0_av_csr.address
		.reset_sequencer_0_av_csr_readdata             (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_readdata),          //  output,   width = 32,                                       .readdata
		.reset_sequencer_0_av_csr_read                 (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_read),              //   input,    width = 1,                                       .read
		.reset_sequencer_0_av_csr_writedata            (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_writedata),         //   input,   width = 32,                                       .writedata
		.reset_sequencer_0_av_csr_write                (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_write),             //   input,    width = 1,                                       .write
		.reset_sequencer_0_av_csr_irq_irq              (),                                                                              //  output,    width = 1,           reset_sequencer_0_av_csr_irq.irq
		.systemclk_f_refclk_fgt_in_refclk_fgt_0        (j204c_f_rx_tx_ip_systemclk_f_refclk_fgt_in_refclk_fgt_0)                        //   input,    width = 1,                 systemclk_f_refclk_fgt.in_refclk_fgt_0
	);

	subsys_jtg_mst jtg_mst (
		.fpga_m_master_address          (jtg_mst_fpga_m_master_address),                            //  output,   width = 32,    fpga_m_master.address
		.fpga_m_master_readdata         (jtg_mst_fpga_m_master_readdata),                           //   input,   width = 32,                 .readdata
		.fpga_m_master_read             (jtg_mst_fpga_m_master_read),                               //  output,    width = 1,                 .read
		.fpga_m_master_write            (jtg_mst_fpga_m_master_write),                              //  output,    width = 1,                 .write
		.fpga_m_master_writedata        (jtg_mst_fpga_m_master_writedata),                          //  output,   width = 32,                 .writedata
		.fpga_m_master_waitrequest      (jtg_mst_fpga_m_master_waitrequest),                        //   input,    width = 1,                 .waitrequest
		.fpga_m_master_readdatavalid    (jtg_mst_fpga_m_master_readdatavalid),                      //   input,    width = 1,                 .readdatavalid
		.fpga_m_master_byteenable       (jtg_mst_fpga_m_master_byteenable),                         //  output,    width = 4,                 .byteenable
		.fpga_m2ocm_pb_s0_waitrequest   (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_waitrequest),   //  output,    width = 1, fpga_m2ocm_pb_s0.waitrequest
		.fpga_m2ocm_pb_s0_readdata      (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_readdata),      //  output,  width = 128,                 .readdata
		.fpga_m2ocm_pb_s0_readdatavalid (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_readdatavalid), //  output,    width = 1,                 .readdatavalid
		.fpga_m2ocm_pb_s0_burstcount    (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_burstcount),    //   input,    width = 1,                 .burstcount
		.fpga_m2ocm_pb_s0_writedata     (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_writedata),     //   input,  width = 128,                 .writedata
		.fpga_m2ocm_pb_s0_address       (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_address),       //   input,   width = 18,                 .address
		.fpga_m2ocm_pb_s0_write         (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_write),         //   input,    width = 1,                 .write
		.fpga_m2ocm_pb_s0_read          (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_read),          //   input,    width = 1,                 .read
		.fpga_m2ocm_pb_s0_byteenable    (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_byteenable),    //   input,   width = 16,                 .byteenable
		.fpga_m2ocm_pb_s0_debugaccess   (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_debugaccess),   //   input,    width = 1,                 .debugaccess
		.fpga_m2ocm_pb_m0_waitrequest   (jtg_mst_fpga_m2ocm_pb_m0_waitrequest),                     //   input,    width = 1, fpga_m2ocm_pb_m0.waitrequest
		.fpga_m2ocm_pb_m0_readdata      (jtg_mst_fpga_m2ocm_pb_m0_readdata),                        //   input,  width = 128,                 .readdata
		.fpga_m2ocm_pb_m0_readdatavalid (jtg_mst_fpga_m2ocm_pb_m0_readdatavalid),                   //   input,    width = 1,                 .readdatavalid
		.fpga_m2ocm_pb_m0_burstcount    (jtg_mst_fpga_m2ocm_pb_m0_burstcount),                      //  output,    width = 1,                 .burstcount
		.fpga_m2ocm_pb_m0_writedata     (jtg_mst_fpga_m2ocm_pb_m0_writedata),                       //  output,  width = 128,                 .writedata
		.fpga_m2ocm_pb_m0_address       (jtg_mst_fpga_m2ocm_pb_m0_address),                         //  output,   width = 18,                 .address
		.fpga_m2ocm_pb_m0_write         (jtg_mst_fpga_m2ocm_pb_m0_write),                           //  output,    width = 1,                 .write
		.fpga_m2ocm_pb_m0_read          (jtg_mst_fpga_m2ocm_pb_m0_read),                            //  output,    width = 1,                 .read
		.fpga_m2ocm_pb_m0_byteenable    (jtg_mst_fpga_m2ocm_pb_m0_byteenable),                      //  output,   width = 16,                 .byteenable
		.fpga_m2ocm_pb_m0_debugaccess   (jtg_mst_fpga_m2ocm_pb_m0_debugaccess),                     //  output,    width = 1,                 .debugaccess
		.hps_m_master_address           (jtg_mst_hps_m_master_address),                             //  output,   width = 32,     hps_m_master.address
		.hps_m_master_readdata          (jtg_mst_hps_m_master_readdata),                            //   input,   width = 32,                 .readdata
		.hps_m_master_read              (jtg_mst_hps_m_master_read),                                //  output,    width = 1,                 .read
		.hps_m_master_write             (jtg_mst_hps_m_master_write),                               //  output,    width = 1,                 .write
		.hps_m_master_writedata         (jtg_mst_hps_m_master_writedata),                           //  output,   width = 32,                 .writedata
		.hps_m_master_waitrequest       (jtg_mst_hps_m_master_waitrequest),                         //   input,    width = 1,                 .waitrequest
		.hps_m_master_readdatavalid     (jtg_mst_hps_m_master_readdatavalid),                       //   input,    width = 1,                 .readdatavalid
		.hps_m_master_byteenable        (jtg_mst_hps_m_master_byteenable),                          //  output,    width = 4,                 .byteenable
		.clk_clk                        (sys_manager_clk_100_out_clk_clk),                          //   input,    width = 1,              clk.clk
		.reset_reset_n                  (~rst_controller_002_reset_out_reset)                       //   input,    width = 1,            reset.reset_n
	);

	subsys_periph periph (
		.ILC_irq_irq                           (periph_ilc_irq_irq),                                 //   input,   width = 2,                        ILC_irq.irq
		.button_pio_external_connection_export (button_pio_external_connection_export),              //   input,   width = 4, button_pio_external_connection.export
		.button_pio_irq_irq                    (irq_mapper_receiver0_irq),                           //  output,   width = 1,                 button_pio_irq.irq
		.dipsw_pio_external_connection_export  (dipsw_pio_external_connection_export),               //   input,   width = 4,  dipsw_pio_external_connection.export
		.dipsw_pio_irq_irq                     (irq_mapper_receiver1_irq),                           //  output,   width = 1,                  dipsw_pio_irq.irq
		.led_pio_external_connection_in_port   (led_pio_external_connection_in_port),                //   input,   width = 3,    led_pio_external_connection.in_port
		.led_pio_external_connection_out_port  (led_pio_external_connection_out_port),               //  output,   width = 3,                               .out_port
		.pb_cpu_0_s0_waitrequest               (mm_interconnect_1_periph_pb_cpu_0_s0_waitrequest),   //  output,   width = 1,                    pb_cpu_0_s0.waitrequest
		.pb_cpu_0_s0_readdata                  (mm_interconnect_1_periph_pb_cpu_0_s0_readdata),      //  output,  width = 32,                               .readdata
		.pb_cpu_0_s0_readdatavalid             (mm_interconnect_1_periph_pb_cpu_0_s0_readdatavalid), //  output,   width = 1,                               .readdatavalid
		.pb_cpu_0_s0_burstcount                (mm_interconnect_1_periph_pb_cpu_0_s0_burstcount),    //   input,   width = 1,                               .burstcount
		.pb_cpu_0_s0_writedata                 (mm_interconnect_1_periph_pb_cpu_0_s0_writedata),     //   input,  width = 32,                               .writedata
		.pb_cpu_0_s0_address                   (mm_interconnect_1_periph_pb_cpu_0_s0_address),       //   input,   width = 9,                               .address
		.pb_cpu_0_s0_write                     (mm_interconnect_1_periph_pb_cpu_0_s0_write),         //   input,   width = 1,                               .write
		.pb_cpu_0_s0_read                      (mm_interconnect_1_periph_pb_cpu_0_s0_read),          //   input,   width = 1,                               .read
		.pb_cpu_0_s0_byteenable                (mm_interconnect_1_periph_pb_cpu_0_s0_byteenable),    //   input,   width = 4,                               .byteenable
		.pb_cpu_0_s0_debugaccess               (mm_interconnect_1_periph_pb_cpu_0_s0_debugaccess),   //   input,   width = 1,                               .debugaccess
		.clk_clk                               (sys_manager_clk_100_out_clk_clk),                    //   input,   width = 1,                            clk.clk
		.reset_reset_n                         (~rst_controller_002_reset_out_reset)                 //   input,   width = 1,                          reset.reset_n
	);

	phipps_peak phipps_peak_0 (
		.clock_bridge_csr_in_clk_clk                                      (clk_ss_0_clk_csr_out_clk_clk),                                                          //   input,    width = 1,                                  clock_bridge_csr_in_clk.clk
		.clock_bridge_dsp_in_clk_clk                                      (clk_ss_0_clk_dsp_out_clk_clk),                                                          //   input,    width = 1,                                  clock_bridge_dsp_in_clk.clk
		.clock_bridge_ecpri_rx_in_clk_clk                                 (clk_ss_0_clk_ftile_402_out_clk_clk),                                                    //   input,    width = 1,                             clock_bridge_ecpri_rx_in_clk.clk
		.clock_bridge_ecpri_tx_in_clk_clk                                 (clk_ss_0_clk_ftile_402_out_clk_clk),                                                    //   input,    width = 1,                             clock_bridge_ecpri_tx_in_clk.clk
		.clock_bridge_eth_in_clk_clk                                      (clk_ss_0_clk_eth_out_clk_clk),                                                          //   input,    width = 1,                                  clock_bridge_eth_in_clk.clk
		.h2f_bridge_s0_waitrequest                                        (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_waitrequest),                             //  output,    width = 1,                                            h2f_bridge_s0.waitrequest
		.h2f_bridge_s0_readdata                                           (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_readdata),                                //  output,   width = 32,                                                         .readdata
		.h2f_bridge_s0_readdatavalid                                      (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_readdatavalid),                           //  output,    width = 1,                                                         .readdatavalid
		.h2f_bridge_s0_burstcount                                         (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_burstcount),                              //   input,    width = 1,                                                         .burstcount
		.h2f_bridge_s0_writedata                                          (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_writedata),                               //   input,   width = 32,                                                         .writedata
		.h2f_bridge_s0_address                                            (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_address),                                 //   input,   width = 23,                                                         .address
		.h2f_bridge_s0_write                                              (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_write),                                   //   input,    width = 1,                                                         .write
		.h2f_bridge_s0_read                                               (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_read),                                    //   input,    width = 1,                                                         .read
		.h2f_bridge_s0_byteenable                                         (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_byteenable),                              //   input,    width = 4,                                                         .byteenable
		.h2f_bridge_s0_debugaccess                                        (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_debugaccess),                             //   input,    width = 1,                                                         .debugaccess
		.h2f_lw_bridge_s0_waitrequest                                     (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_waitrequest),                          //  output,    width = 1,                                         h2f_lw_bridge_s0.waitrequest
		.h2f_lw_bridge_s0_readdata                                        (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_readdata),                             //  output,   width = 32,                                                         .readdata
		.h2f_lw_bridge_s0_readdatavalid                                   (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_readdatavalid),                        //  output,    width = 1,                                                         .readdatavalid
		.h2f_lw_bridge_s0_burstcount                                      (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_burstcount),                           //   input,    width = 1,                                                         .burstcount
		.h2f_lw_bridge_s0_writedata                                       (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_writedata),                            //   input,   width = 32,                                                         .writedata
		.h2f_lw_bridge_s0_address                                         (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_address),                              //   input,   width = 20,                                                         .address
		.h2f_lw_bridge_s0_write                                           (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_write),                                //   input,    width = 1,                                                         .write
		.h2f_lw_bridge_s0_read                                            (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_read),                                 //   input,    width = 1,                                                         .read
		.h2f_lw_bridge_s0_byteenable                                      (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_byteenable),                           //   input,    width = 4,                                                         .byteenable
		.h2f_lw_bridge_s0_debugaccess                                     (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_debugaccess),                          //   input,    width = 1,                                                         .debugaccess
		.csr_in_reset_reset_n                                             (rst_ss_0_rst_csr_out_reset_reset),                                                      //   input,    width = 1,                                             csr_in_reset.reset_n
		.dsp_in_reset_reset_n                                             (~rst_ss_0_dsp_rst_cntrl_reset_out_reset),                                               //   input,    width = 1,                                             dsp_in_reset.reset_n
		.eth_in_reset_reset_n                                             (~rst_ss_0_eth_rst_cntrl_reset_out_reset),                                               //   input,    width = 1,                                             eth_in_reset.reset_n
		.rst_ecpri_n_reset_n                                              (~rst_ss_0_ecpri_rst_cntrl_reset_out_reset),                                             //   input,    width = 1,                                              rst_ecpri_n.reset_n
		.radio_config_status_dup2_radio_config_status                     (phipps_peak_0_radio_config_status_dup2_radio_config_status),                            //  output,   width = 56,                                 radio_config_status_dup2.radio_config_status
		.rst_soft_n_dup4_rst_soft_n                                       (phipps_peak_0_rst_soft_n_dup4_rst_soft_n),                                              //  output,    width = 1,                                          rst_soft_n_dup4.rst_soft_n
		.interface_sel_data                                               (dfd_subsystem_interface_sel_data),                                                      //   input,   width = 32,                                            interface_sel.data
		.ddc_avst_sink_avst_sink_valid                                    (ddc_avst_sink_avst_sink_valid),                                                         //   input,    width = 1,                                            ddc_avst_sink.avst_sink_valid
		.ddc_avst_sink_avst_sink_channel                                  (ddc_avst_sink_avst_sink_channel),                                                       //   input,    width = 8,                                                         .avst_sink_channel
		.ddc_avst_sink_avst_sink_data_l1                                  (ddc_avst_sink_avst_sink_data_l1),                                                       //   input,   width = 32,                                                         .avst_sink_data_l1
		.ddc_avst_sink_avst_sink_data_l2                                  (ddc_avst_sink_avst_sink_data_l2),                                                       //   input,   width = 32,                                                         .avst_sink_data_l2
		.ddc_avst_sink_avst_sink_data_l3                                  (ddc_avst_sink_avst_sink_data_l3),                                                       //   input,   width = 32,                                                         .avst_sink_data_l3
		.ddc_avst_sink_avst_sink_data_l4                                  (ddc_avst_sink_avst_sink_data_l4),                                                       //   input,   width = 32,                                                         .avst_sink_data_l4
		.ddc_avst_sink_avst_sink_data_l5                                  (ddc_avst_sink_avst_sink_data_l5),                                                       //   input,   width = 32,                                                         .avst_sink_data_l5
		.ddc_avst_sink_avst_sink_data_l6                                  (ddc_avst_sink_avst_sink_data_l6),                                                       //   input,   width = 32,                                                         .avst_sink_data_l6
		.ddc_avst_sink_avst_sink_data_l7                                  (ddc_avst_sink_avst_sink_data_l7),                                                       //   input,   width = 32,                                                         .avst_sink_data_l7
		.ddc_avst_sink_avst_sink_data_l8                                  (ddc_avst_sink_avst_sink_data_l8),                                                       //   input,   width = 32,                                                         .avst_sink_data_l8
		.duc_avst_source_duc_avst_source_valid                            (duc_avst_source_duc_avst_source_valid),                                                 //  output,    width = 1,                                          duc_avst_source.duc_avst_source_valid
		.duc_avst_source_duc_avst_source_data0                            (duc_avst_source_duc_avst_source_data0),                                                 //  output,   width = 32,                                                         .duc_avst_source_data0
		.duc_avst_source_duc_avst_source_data1                            (duc_avst_source_duc_avst_source_data1),                                                 //  output,   width = 32,                                                         .duc_avst_source_data1
		.duc_avst_source_duc_avst_source_data2                            (duc_avst_source_duc_avst_source_data2),                                                 //  output,   width = 32,                                                         .duc_avst_source_data2
		.duc_avst_source_duc_avst_source_data3                            (duc_avst_source_duc_avst_source_data3),                                                 //  output,   width = 32,                                                         .duc_avst_source_data3
		.duc_avst_source_duc_avst_source_data4                            (duc_avst_source_duc_avst_source_data4),                                                 //  output,   width = 32,                                                         .duc_avst_source_data4
		.duc_avst_source_duc_avst_source_data5                            (duc_avst_source_duc_avst_source_data5),                                                 //  output,   width = 32,                                                         .duc_avst_source_data5
		.duc_avst_source_duc_avst_source_data6                            (duc_avst_source_duc_avst_source_data6),                                                 //  output,   width = 32,                                                         .duc_avst_source_data6
		.duc_avst_source_duc_avst_source_data7                            (duc_avst_source_duc_avst_source_data7),                                                 //  output,   width = 32,                                                         .duc_avst_source_data7
		.duc_avst_source_duc_avst_source_channel                          (duc_avst_source_duc_avst_source_channel),                                               //  output,    width = 8,                                                         .duc_avst_source_channel
		.dxc_ss_top_0_rfp_pulse_data                                      (tod_subsys_0_tod_timestamp_96b_0_rfp_sync_pul_data),                                    //   input,    width = 1,                                   dxc_ss_top_0_rfp_pulse.data
		.dxc_avst_selctd_cap_intf_valid                                   (phipps_peak_0_dxc_avst_selctd_cap_intf_valid),                                          //  output,    width = 1,                                 dxc_avst_selctd_cap_intf.valid
		.dxc_avst_selctd_cap_intf_data                                    (phipps_peak_0_dxc_avst_selctd_cap_intf_data),                                           //  output,   width = 32,                                                         .data
		.dxc_avst_selctd_cap_intf_channel                                 (phipps_peak_0_dxc_avst_selctd_cap_intf_channel),                                        //  output,    width = 3,                                                         .channel
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_skip_crc              (avst_tx_ptp_i_av_st_tx_skip_crc),                                                       //   input,    width = 1,                          avst_axist_bridge_0_avst_tx_ptp.i_av_st_tx_skip_crc
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_ts_valid          (avst_tx_ptp_i_av_st_tx_ptp_ts_valid),                                                   //   input,    width = 2,                                                         .i_av_st_tx_ptp_ts_valid
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_ins_ets           (avst_tx_ptp_i_av_st_tx_ptp_ins_ets),                                                    //   input,    width = 1,                                                         .i_av_st_tx_ptp_ins_ets
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_ins_cf            (avst_tx_ptp_i_av_st_tx_ptp_ins_cf),                                                     //   input,    width = 1,                                                         .i_av_st_tx_ptp_ins_cf
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_tx_its            (avst_tx_ptp_i_av_st_tx_ptp_tx_its),                                                     //   input,   width = 96,                                                         .i_av_st_tx_ptp_tx_its
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_asym_p2p_idx      (avst_tx_ptp_i_av_st_tx_ptp_asym_p2p_idx),                                               //   input,    width = 7,                                                         .i_av_st_tx_ptp_asym_p2p_idx
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_asym_sign         (avst_tx_ptp_i_av_st_tx_ptp_asym_sign),                                                  //   input,    width = 1,                                                         .i_av_st_tx_ptp_asym_sign
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_asym              (avst_tx_ptp_i_av_st_tx_ptp_asym),                                                       //   input,    width = 1,                                                         .i_av_st_tx_ptp_asym
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_p2p               (avst_tx_ptp_i_av_st_tx_ptp_p2p),                                                        //   input,    width = 1,                                                         .i_av_st_tx_ptp_p2p
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_ts_format         (avst_tx_ptp_i_av_st_tx_ptp_ts_format),                                                  //   input,    width = 1,                                                         .i_av_st_tx_ptp_ts_format
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_update_eb         (avst_tx_ptp_i_av_st_tx_ptp_update_eb),                                                  //   input,    width = 1,                                                         .i_av_st_tx_ptp_update_eb
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_zero_csum         (avst_tx_ptp_i_av_st_tx_ptp_zero_csum),                                                  //   input,    width = 1,                                                         .i_av_st_tx_ptp_zero_csum
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_eb_offset         (avst_tx_ptp_i_av_st_tx_ptp_eb_offset),                                                  //   input,   width = 16,                                                         .i_av_st_tx_ptp_eb_offset
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_csum_offset       (avst_tx_ptp_i_av_st_tx_ptp_csum_offset),                                                //   input,   width = 16,                                                         .i_av_st_tx_ptp_csum_offset
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_cf_offset         (avst_tx_ptp_i_av_st_tx_ptp_cf_offset),                                                  //   input,   width = 16,                                                         .i_av_st_tx_ptp_cf_offset
		.avst_axist_bridge_0_avst_tx_ptp_i_av_st_tx_ptp_ts_offset         (avst_tx_ptp_i_av_st_tx_ptp_ts_offset),                                                  //   input,   width = 16,                                                         .i_av_st_tx_ptp_ts_offset
		.avst_axist_bridge_0_axit_tx_if_tready                            (avst_axist_bridge_0_axit_tx_if_tready),                                                 //   input,    width = 1,                           avst_axist_bridge_0_axit_tx_if.tready
		.avst_axist_bridge_0_axit_tx_if_tvalid                            (avst_axist_bridge_0_axit_tx_if_tvalid),                                                 //  output,    width = 1,                                                         .tvalid
		.avst_axist_bridge_0_axit_tx_if_tdata                             (avst_axist_bridge_0_axit_tx_if_tdata),                                                  //  output,   width = 64,                                                         .tdata
		.avst_axist_bridge_0_axit_tx_if_tlast                             (avst_axist_bridge_0_axit_tx_if_tlast),                                                  //  output,    width = 1,                                                         .tlast
		.avst_axist_bridge_0_axit_tx_if_tkeep                             (avst_axist_bridge_0_axit_tx_if_tkeep),                                                  //  output,    width = 8,                                                         .tkeep
		.avst_axist_bridge_0_axit_tx_if_tuser                             (avst_axist_bridge_0_axit_tx_if_tuser),                                                  //  output,    width = 2,                                                         .tuser
		.avst_axist_bridge_0_axist_tx_user_o_axi_st_tx_tuser_ptp          (axist_tx_user_o_axi_st_tx_tuser_ptp),                                                   //  output,   width = 94,                        avst_axist_bridge_0_axist_tx_user.o_axi_st_tx_tuser_ptp
		.avst_axist_bridge_0_axist_tx_user_o_axi_st_tx_tuser_ptp_extended (axist_tx_user_o_axi_st_tx_tuser_ptp_extended),                                          //  output,  width = 328,                                                         .o_axi_st_tx_tuser_ptp_extended
		.avst_axist_bridge_0_avst_rx_ptp_o_av_st_rxstatus_data            (avst_rx_ptp_o_av_st_rxstatus_data),                                                     //  output,   width = 40,                          avst_axist_bridge_0_avst_rx_ptp.o_av_st_rxstatus_data
		.avst_axist_bridge_0_avst_rx_ptp_o_av_st_rxstatus_valid           (avst_rx_ptp_o_av_st_rxstatus_valid),                                                    //  output,    width = 1,                                                         .o_av_st_rxstatus_valid
		.avst_axist_bridge_0_avst_rx_ptp_o_av_st_ptp_rx_its               (avst_rx_ptp_o_av_st_ptp_rx_its),                                                        //  output,   width = 96,                                                         .o_av_st_ptp_rx_its
		.avst_axist_bridge_0_axist_rx_if_tvalid                           (hssi_ss_1_p0_axi_st_rx_interface_tvalid),                                               //   input,    width = 1,                          avst_axist_bridge_0_axist_rx_if.tvalid
		.avst_axist_bridge_0_axist_rx_if_tdata                            (hssi_ss_1_p0_axi_st_rx_interface_tdata),                                                //   input,   width = 64,                                                         .tdata
		.avst_axist_bridge_0_axist_rx_if_tlast                            (hssi_ss_1_p0_axi_st_rx_interface_tlast),                                                //   input,    width = 1,                                                         .tlast
		.avst_axist_bridge_0_axist_rx_if_tkeep                            (hssi_ss_1_p0_axi_st_rx_interface_tkeep),                                                //   input,    width = 8,                                                         .tkeep
		.avst_axist_bridge_0_axist_rx_if_tuser                            (hssi_ss_1_p0_axi_st_rx_interface_tuser),                                                //   input,    width = 7,                                                         .tuser
		.avst_axist_bridge_0_axist_rx_user_i_axi_st_rx_tuser_sts          (axist_rx_user_i_axi_st_rx_tuser_sts),                                                   //   input,    width = 5,                        avst_axist_bridge_0_axist_rx_user.i_axi_st_rx_tuser_sts
		.avst_axist_bridge_0_axist_rx_user_i_axi_st_rx_tuser_sts_extended (axist_rx_user_i_axi_st_rx_tuser_sts_extended),                                          //   input,   width = 32,                                                         .i_axi_st_rx_tuser_sts_extended
		.avst_axist_bridge_0_axist_rx_user_i_axi_st_rx_ingrts0_tdata      (axist_rx_user_i_axi_st_rx_ingrts0_tdata),                                               //   input,   width = 96,                                                         .i_axi_st_rx_ingrts0_tdata
		.avst_axist_bridge_0_axist_rx_user_i_axi_st_rx_ingrts0_tvalid     (axist_rx_user_i_axi_st_rx_ingrts0_tvalid),                                              //   input,    width = 1,                                                         .i_axi_st_rx_ingrts0_tvalid
		.ecpri_ext_sink_valid                                             (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid),         //   input,    width = 1,                                           ecpri_ext_sink.valid
		.ecpri_ext_sink_data                                              (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data),          //   input,   width = 64,                                                         .data
		.ecpri_ext_sink_startofpacket                                     (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket), //   input,    width = 1,                                                         .startofpacket
		.ecpri_ext_sink_endofpacket                                       (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket),   //   input,    width = 1,                                                         .endofpacket
		.ecpri_ext_sink_empty                                             (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty),         //   input,    width = 3,                                                         .empty
		.ecpri_ext_sink_error                                             (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error),         //   input,    width = 1,                                                         .error
		.ecpri_ext_sink_ready                                             (dma_subsys_dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready),         //  output,    width = 1,                                                         .ready
		.ecpri_ext_source_valid                                           (phipps_peak_0_ecpri_ext_source_valid),                                                  //  output,    width = 1,                                         ecpri_ext_source.valid
		.ecpri_ext_source_data                                            (phipps_peak_0_ecpri_ext_source_data),                                                   //  output,   width = 64,                                                         .data
		.ecpri_ext_source_startofpacket                                   (phipps_peak_0_ecpri_ext_source_startofpacket),                                          //  output,    width = 1,                                                         .startofpacket
		.ecpri_ext_source_endofpacket                                     (phipps_peak_0_ecpri_ext_source_endofpacket),                                            //  output,    width = 1,                                                         .endofpacket
		.ecpri_ext_source_empty                                           (phipps_peak_0_ecpri_ext_source_empty),                                                  //  output,    width = 3,                                                         .empty
		.ecpri_ext_source_error                                           (phipps_peak_0_ecpri_ext_source_error),                                                  //  output,    width = 6,                                                         .error
		.ptp_tod_concat_out_o_mac_ptp_fp                                  (ptp_tod_concat_out_o_mac_ptp_fp),                                                       //  output,   width = 22,                                       ptp_tod_concat_out.o_mac_ptp_fp
		.ptp_tod_concat_out_o_mac_ptp_ts_req                              (ptp_tod_concat_out_o_mac_ptp_ts_req),                                                   //  output,    width = 1,                                                         .o_mac_ptp_ts_req
		.ptp_tod_concat_out_i_mac_ptp_tx_ets_valid                        (ptp_tod_concat_out_i_mac_ptp_tx_ets_valid),                                             //   input,    width = 1,                                                         .i_mac_ptp_tx_ets_valid
		.ptp_tod_concat_out_i_mac_ptp_tx_ets                              (ptp_tod_concat_out_i_mac_ptp_tx_ets),                                                   //   input,   width = 96,                                                         .i_mac_ptp_tx_ets
		.ptp_tod_concat_out_i_mac_ptp_tx_ets_fp                           (ptp_tod_concat_out_i_mac_ptp_tx_ets_fp),                                                //   input,   width = 22,                                                         .i_mac_ptp_tx_ets_fp
		.ptp_tod_concat_out_i_mac_ptp_rx_its_valid                        (ptp_tod_concat_out_i_mac_ptp_rx_its_valid),                                             //   input,    width = 1,                                                         .i_mac_ptp_rx_its_valid
		.ptp_tod_concat_out_i_mac_ptp_rx_its                              (ptp_tod_concat_out_i_mac_ptp_rx_its),                                                   //   input,   width = 96,                                                         .i_mac_ptp_rx_its
		.ptp_tod_concat_out_i_ext_ptp_fp                                  (ptp_tod_concat_out_i_ext_ptp_fp),                                                       //   input,   width = 20,                                                         .i_ext_ptp_fp
		.ptp_tod_concat_out_i_ext_ptp_ts_req                              (ptp_tod_concat_out_i_ext_ptp_ts_req),                                                   //   input,    width = 1,                                                         .i_ext_ptp_ts_req
		.ptp_tod_concat_out_o_ext_ptp_tx_ets_valid                        (ptp_tod_concat_out_o_ext_ptp_tx_ets_valid),                                             //  output,    width = 1,                                                         .o_ext_ptp_tx_ets_valid
		.ptp_tod_concat_out_o_ext_ptp_tx_ets                              (ptp_tod_concat_out_o_ext_ptp_tx_ets),                                                   //  output,   width = 96,                                                         .o_ext_ptp_tx_ets
		.ptp_tod_concat_out_o_ext_ptp_tx_ets_fp                           (ptp_tod_concat_out_o_ext_ptp_tx_ets_fp),                                                //  output,   width = 20,                                                         .o_ext_ptp_tx_ets_fp
		.ptp_tod_concat_out_o_ext_ptp_rx_its                              (ptp_tod_concat_out_o_ext_ptp_rx_its),                                                   //  output,   width = 96,                                                         .o_ext_ptp_rx_its
		.ptp_tod_concat_out_o_ext_ptp_rx_its_valid                        (ptp_tod_concat_out_o_ext_ptp_rx_its_valid),                                             //  output,    width = 1,                                                         .o_ext_ptp_rx_its_valid
		.rx_pcs_ready_rx_pcs_ready                                        (phipps_peak_0_rx_pcs_ready_rx_pcs_ready),                                               //   input,    width = 1,                                             rx_pcs_ready.rx_pcs_ready
		.tx_lanes_stable_tx_lanes_stable                                  (phipps_peak_0_tx_lanes_stable_tx_lanes_stable),                                         //   input,    width = 1,                                          tx_lanes_stable.tx_lanes_stable
		.ecpri_oran_top_0_oran_tx_tod_96b_data_tdata                      (tod_subsys_0_tx_oran_tod_time_of_day_96b_tdata),                                        //   input,   width = 96,                    ecpri_oran_top_0_oran_tx_tod_96b_data.tdata
		.ecpri_oran_top_0_oran_tx_tod_96b_data_tvalid                     (tod_subsys_0_tx_oran_tod_time_of_day_96b_tvalid),                                       //   input,    width = 1,                                                         .tvalid
		.ecpri_oran_top_0_oran_rx_tod_96b_data_tdata                      (tod_subsys_0_rx_oran_tod_time_of_day_96b_tdata),                                        //   input,   width = 96,                    ecpri_oran_top_0_oran_rx_tod_96b_data.tdata
		.ecpri_oran_top_0_oran_rx_tod_96b_data_tvalid                     (tod_subsys_0_rx_oran_tod_time_of_day_96b_tvalid),                                       //   input,    width = 1,                                                         .tvalid
		.xran_timestamp_tod_in_data                                       (tod_subsys_0_cdc_pipeline_0_dataout_data),                                              //   input,   width = 96,                                    xran_timestamp_tod_in.data
		.timeout_cntr_intr_uplane_irq                                     (irq_mapper_receiver13_irq),                                                             //  output,    width = 1,                                 timeout_cntr_intr_uplane.irq
		.timeout_cntr_intr_cplane_irq                                     (irq_mapper_receiver12_irq),                                                             //  output,    width = 1,                                 timeout_cntr_intr_cplane.irq
		.fifo_full_intr_irq                                               (irq_mapper_receiver4_irq),                                                              //  output,    width = 1,                                           fifo_full_intr.irq
		.pwr_mtr_h2f_bridge_s0_waitrequest                                (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_waitrequest),                     //  output,    width = 1,                                    pwr_mtr_h2f_bridge_s0.waitrequest
		.pwr_mtr_h2f_bridge_s0_readdata                                   (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdata),                        //  output,   width = 32,                                                         .readdata
		.pwr_mtr_h2f_bridge_s0_readdatavalid                              (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdatavalid),                   //  output,    width = 1,                                                         .readdatavalid
		.pwr_mtr_h2f_bridge_s0_burstcount                                 (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_burstcount),                      //   input,    width = 1,                                                         .burstcount
		.pwr_mtr_h2f_bridge_s0_writedata                                  (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_writedata),                       //   input,   width = 32,                                                         .writedata
		.pwr_mtr_h2f_bridge_s0_address                                    (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_address),                         //   input,   width = 17,                                                         .address
		.pwr_mtr_h2f_bridge_s0_write                                      (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_write),                           //   input,    width = 1,                                                         .write
		.pwr_mtr_h2f_bridge_s0_read                                       (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_read),                            //   input,    width = 1,                                                         .read
		.pwr_mtr_h2f_bridge_s0_byteenable                                 (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_byteenable),                      //   input,    width = 4,                                                         .byteenable
		.pwr_mtr_h2f_bridge_s0_debugaccess                                (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_debugaccess),                     //   input,    width = 1,                                                         .debugaccess
		.lphy_ss_top_0_pb_avst_sink_valid                                 (),                                                                                      //   input,    width = 1,                               lphy_ss_top_0_pb_avst_sink.valid
		.lphy_ss_top_0_pb_avst_sink_data                                  (),                                                                                      //   input,   width = 64,                                                         .data
		.lphy_ss_top_0_pb_avst_sink_ready                                 (),                                                                                      //  output,    width = 1,                                                         .ready
		.lphy_avst_selctd_cap_intf_valid                                  (phipps_peak_0_lphy_avst_selctd_cap_intf_valid),                                         //  output,    width = 1,                                lphy_avst_selctd_cap_intf.valid
		.lphy_avst_selctd_cap_intf_data                                   (phipps_peak_0_lphy_avst_selctd_cap_intf_data),                                          //  output,   width = 32,                                                         .data
		.lphy_avst_selctd_cap_intf_channel                                (phipps_peak_0_lphy_avst_selctd_cap_intf_channel),                                       //  output,    width = 3,                                                         .channel
		.lphy_ss_top_0_frame_status_counter_reset_data                    (tod_subsys_0_tod_timestamp_96b_0_rfp_sync_pul_dup_data),                                //   input,    width = 1,                 lphy_ss_top_0_frame_status_counter_reset.data
		.lphy_ss_top_0_lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l1_irq     (irq_mapper_receiver9_irq),                                                              //  output,    width = 1, lphy_ss_top_0_lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l1.irq
		.lphy_ss_top_0_lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l2_irq     (irq_mapper_receiver10_irq),                                                             //  output,    width = 1, lphy_ss_top_0_lphy_ss_top_pwr_mtr_ifft_hist_done_intr_l2.irq
		.lphy_ss_top_0_lphy_ss_top_pwr_mtr_fft_hist_done_intr_l1_irq      (irq_mapper_receiver7_irq),                                                              //  output,    width = 1,  lphy_ss_top_0_lphy_ss_top_pwr_mtr_fft_hist_done_intr_l1.irq
		.lphy_ss_top_0_lphy_ss_top_pwr_mtr_fft_hist_done_intr_l2_irq      (irq_mapper_receiver8_irq),                                                              //  output,    width = 1,  lphy_ss_top_0_lphy_ss_top_pwr_mtr_fft_hist_done_intr_l2.irq
		.lphy_ss_top_0_lphy_ss_top_duc_ddc_lpbk_en_data                   (phipps_peak_0_lphy_ss_top_0_lphy_ss_top_duc_ddc_lpbk_en_data)                           //  output,    width = 1,                lphy_ss_top_0_lphy_ss_top_duc_ddc_lpbk_en.data
	);

	rst_ss rst_ss_0 (
		.dsp_rst_cntrl_reset_in0_reset         (rst_dsp_in_reset_reset),                   //   input,  width = 1,         dsp_rst_cntrl_reset_in0.reset
		.dsp_rst_cntrl_clk_clk                 (clk_ss_0_clk_dsp_out_clk_clk),             //   input,  width = 1,               dsp_rst_cntrl_clk.clk
		.dsp_rst_cntrl_reset_out_reset         (rst_ss_0_dsp_rst_cntrl_reset_out_reset),   //  output,  width = 1,         dsp_rst_cntrl_reset_out.reset
		.ecpri_rst_cntrl_reset_in0_reset       (~hssi_ss_1_o_p0_ereset_n_reset),           //   input,  width = 1,       ecpri_rst_cntrl_reset_in0.reset
		.ecpri_rst_cntrl_clk_clk               (clk_ss_0_clk_ftile_402_out_clk_clk),       //   input,  width = 1,             ecpri_rst_cntrl_clk.clk
		.ecpri_rst_cntrl_reset_out_reset       (rst_ss_0_ecpri_rst_cntrl_reset_out_reset), //  output,  width = 1,       ecpri_rst_cntrl_reset_out.reset
		.eth_rst_cntrl_reset_in0_reset         (rst_eth_in_reset_reset),                   //   input,  width = 1,         eth_rst_cntrl_reset_in0.reset
		.eth_rst_cntrl_clk_clk                 (clk_ss_0_clk_eth_out_clk_clk),             //   input,  width = 1,               eth_rst_cntrl_clk.clk
		.eth_rst_cntrl_reset_out_reset         (rst_ss_0_eth_rst_cntrl_reset_out_reset),   //  output,  width = 1,         eth_rst_cntrl_reset_out.reset
		.reset_bridge_act_high_clk_clk         (clk_ss_0_clk_csr_out_clk_clk),             //   input,  width = 1,       reset_bridge_act_high_clk.clk
		.reset_bridge_act_high_in_reset_reset  (rst_csr_act_high_in_reset_reset),          //   input,  width = 1,  reset_bridge_act_high_in_reset.reset
		.reset_bridge_act_high_out_reset_reset (),                                         //  output,  width = 1, reset_bridge_act_high_out_reset.reset
		.rst_csr_clk_clk                       (clk_ss_0_clk_csr_out_clk_clk),             //   input,  width = 1,                     rst_csr_clk.clk
		.rst_csr_in_reset_reset_n              (rst_csr_in_reset_reset_n),                 //   input,  width = 1,                rst_csr_in_reset.reset_n
		.rst_csr_out_reset_reset_n             (rst_ss_0_rst_csr_out_reset_reset),         //  output,  width = 1,               rst_csr_out_reset.reset_n
		.reset_bridge_rec_rx_clk_clk           (hssi_ss_1_o_p0_clk_rec_div_clk_signal),    //   input,  width = 1,         reset_bridge_rec_rx_clk.clk
		.reset_bridge_rec_rx_in_reset_reset    (rst_controller_003_reset_out_reset),       //   input,  width = 1,    reset_bridge_rec_rx_in_reset.reset
		.reset_bridge_rec_rx_out_reset_reset   (),                                         //  output,  width = 1,   reset_bridge_rec_rx_out_reset.reset
		.reset_bridge_tx_div_clk_clk           (hssi_ss_1_o_p0_clk_tx_div_clk),            //   input,  width = 1,         reset_bridge_tx_div_clk.clk
		.reset_bridge_tx_div_in_reset_reset    (rst_controller_004_reset_out_reset),       //   input,  width = 1,    reset_bridge_tx_div_in_reset.reset
		.reset_bridge_tx_div_out_reset_reset   ()                                          //  output,  width = 1,   reset_bridge_tx_div_out_reset.reset
	);

	sys_manager sys_manager (
		.clk_100_in_clk_clk                               (clk_100_clk),                                                //   input,   width = 1,                           clk_100_in_clk.clk
		.clk_100_out_clk_clk                              (sys_manager_clk_100_out_clk_clk),                            //  output,   width = 1,                          clk_100_out_clk.clk
		.dma_subsys_port0_rx_dma_resetn_clk_clk           (sys_manager_clk_100_out_clk_clk),                            //   input,   width = 1,       dma_subsys_port0_rx_dma_resetn_clk.clk
		.dma_subsys_port0_rx_dma_resetn_in_reset_reset_n  (dma_subsys_port0_rx_dma_resetn_reset_n),                     //   input,   width = 1,  dma_subsys_port0_rx_dma_resetn_in_reset.reset_n
		.dma_subsys_port0_rx_dma_resetn_out_reset_reset_n (sys_manager_dma_subsys_port0_rx_dma_resetn_out_reset_reset), //  output,   width = 1, dma_subsys_port0_rx_dma_resetn_out_reset.reset_n
		.dma_subsys_port1_rx_dma_resetn_clk_clk           (sys_manager_clk_100_out_clk_clk),                            //   input,   width = 1,       dma_subsys_port1_rx_dma_resetn_clk.clk
		.dma_subsys_port1_rx_dma_resetn_in_reset_reset_n  (dma_subsys_port1_rx_dma_resetn_reset_n),                     //   input,   width = 1,  dma_subsys_port1_rx_dma_resetn_in_reset.reset_n
		.dma_subsys_port1_rx_dma_resetn_out_reset_reset_n (sys_manager_dma_subsys_port1_rx_dma_resetn_out_reset_reset), //  output,   width = 1, dma_subsys_port1_rx_dma_resetn_out_reset.reset_n
		.ftile_iopll_ptp_sampling_refclk_clk              (sys_manager_clk_100_out_clk_clk),                            //   input,   width = 1,          ftile_iopll_ptp_sampling_refclk.clk
		.ftile_iopll_ptp_sampling_reset_reset             (~sys_manager_rst_in_out_reset_reset),                        //   input,   width = 1,           ftile_iopll_ptp_sampling_reset.reset
		.ftile_iopll_ptp_sampling_outclk0_clk             (sys_manager_ftile_iopll_ptp_sampling_outclk0_clk),           //  output,   width = 1,         ftile_iopll_ptp_sampling_outclk0.clk
		.ftile_iopll_todsync_sampling_refclk_clk          (sys_manager_qsys_top_master_todclk_0_out_clk_clk),           //   input,   width = 1,      ftile_iopll_todsync_sampling_refclk.clk
		.ftile_iopll_todsync_sampling_locked_lock         (sys_manager_ftile_iopll_todsync_sampling_locked_lock),       //  output,   width = 1,      ftile_iopll_todsync_sampling_locked.lock
		.ftile_iopll_todsync_sampling_reset_reset         (~sys_manager_rst_in_out_reset_reset),                        //   input,   width = 1,       ftile_iopll_todsync_sampling_reset.reset
		.ftile_iopll_todsync_sampling_outclk0_clk         (sys_manager_ftile_iopll_todsync_sampling_outclk0_clk),       //  output,   width = 1,     ftile_iopll_todsync_sampling_outclk0.clk
		.qsys_top_master_todclk_0_in_clk_clk              (qsys_top_master_todclk_0_in_clk_clk),                        //   input,   width = 1,          qsys_top_master_todclk_0_in_clk.clk
		.qsys_top_master_todclk_0_out_clk_clk             (sys_manager_qsys_top_master_todclk_0_out_clk_clk),           //  output,   width = 1,         qsys_top_master_todclk_0_out_clk.clk
		.rst_in_clk_clk                                   (sys_manager_clk_100_out_clk_clk),                            //   input,   width = 1,                               rst_in_clk.clk
		.rst_in_in_reset_reset_n                          (reset_reset_n),                                              //   input,   width = 1,                          rst_in_in_reset.reset_n
		.rst_in_out_reset_reset_n                         (sys_manager_rst_in_out_reset_reset),                         //  output,   width = 1,                         rst_in_out_reset.reset_n
		.sysid_clk_clk                                    (sys_manager_clk_100_out_clk_clk),                            //   input,   width = 1,                                sysid_clk.clk
		.sysid_reset_reset_n                              (~rst_controller_reset_out_reset),                            //   input,   width = 1,                              sysid_reset.reset_n
		.sysid_control_slave_readdata                     (mm_interconnect_1_sys_manager_sysid_control_slave_readdata), //  output,  width = 32,                      sysid_control_slave.readdata
		.sysid_control_slave_address                      (mm_interconnect_1_sys_manager_sysid_control_slave_address),  //   input,   width = 1,                                         .address
		.user_rst_clkgate_0_ninit_done_ninit_done         (ninit_done_ninit_done)                                       //  output,   width = 1,            user_rst_clkgate_0_ninit_done.ninit_done
	);

	tod_subsys tod_subsys_0 (
		.cdc_pipeline_0_dst_clk_clk                              (clk_ss_0_clk_ftile_402_out_clk_clk),                                                     //   input,   width = 1,                             cdc_pipeline_0_dst_clk.clk
		.cdc_pipeline_0_rst_dst_clk_n_reset_n                    (~rst_ss_0_eth_rst_cntrl_reset_out_reset),                                                //   input,   width = 1,                       cdc_pipeline_0_rst_dst_clk_n.reset_n
		.cdc_pipeline_0_dataout_data                             (tod_subsys_0_cdc_pipeline_0_dataout_data),                                               //  output,  width = 96,                             cdc_pipeline_0_dataout.data
		.clock_bridge_100_in_clk_clk                             (clk_ss_0_clk_csr_out_clk_clk),                                                           //   input,   width = 1,                            clock_bridge_100_in_clk.clk
		.clock_bridge_156_in_clk_clk                             (sys_manager_qsys_top_master_todclk_0_out_clk_clk),                                       //   input,   width = 1,                            clock_bridge_156_in_clk.clk
		.reset_bridge_100_in_reset_reset_n                       (rst_ss_0_rst_csr_out_reset_reset),                                                       //   input,   width = 1,                          reset_bridge_100_in_reset.reset_n
		.reset_bridge_156_in_reset_reset                         (rst_controller_005_reset_out_reset),                                                     //   input,   width = 1,                          reset_bridge_156_in_reset.reset
		.tod_timestamp_96b_0_pps_in_pps_in                       (tod_timestamp_96b_0_pps_in_pps_in),                                                      //   input,   width = 1,                         tod_timestamp_96b_0_pps_in.pps_in
		.tod_timestamp_96b_0_rfp_sync_pul_data                   (tod_subsys_0_tod_timestamp_96b_0_rfp_sync_pul_data),                                     //  output,   width = 1,                   tod_timestamp_96b_0_rfp_sync_pul.data
		.tod_timestamp_96b_0_tod_timestamp_96b_csr_address       (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_address),       //   input,   width = 5,          tod_timestamp_96b_0_tod_timestamp_96b_csr.address
		.tod_timestamp_96b_0_tod_timestamp_96b_csr_write         (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_write),         //   input,   width = 1,                                                   .write
		.tod_timestamp_96b_0_tod_timestamp_96b_csr_read          (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_read),          //   input,   width = 1,                                                   .read
		.tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata     (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata),     //   input,  width = 32,                                                   .writedata
		.tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata      (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata),      //  output,  width = 32,                                                   .readdata
		.tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest   (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest),   //  output,   width = 1,                                                   .waitrequest
		.tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid), //  output,   width = 1,                                                   .readdatavalid
		.tod_timestamp_96b_0_rfp_sync_pul_dup_data               (tod_subsys_0_tod_timestamp_96b_0_rfp_sync_pul_dup_data),                                 //  output,   width = 1,               tod_timestamp_96b_0_rfp_sync_pul_dup.data
		.master_tod_top_0_csr_write                              (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_write),                              //   input,   width = 1,                               master_tod_top_0_csr.write
		.master_tod_top_0_csr_writedata                          (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_writedata),                          //   input,  width = 32,                                                   .writedata
		.master_tod_top_0_csr_read                               (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_read),                               //   input,   width = 1,                                                   .read
		.master_tod_top_0_csr_readdata                           (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_readdata),                           //  output,  width = 32,                                                   .readdata
		.master_tod_top_0_csr_waitrequest                        (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_waitrequest),                        //  output,   width = 1,                                                   .waitrequest
		.master_tod_top_0_csr_address                            (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_address),                            //   input,   width = 4,                                                   .address
		.master_tod_top_0_i_reconfig_rst_n_reset_n               (~rst_controller_002_reset_out_reset),                                                    //   input,   width = 1,                  master_tod_top_0_i_reconfig_rst_n.reset_n
		.master_tod_top_0_pulse_per_second_pps                   (master_tod_top_0_pulse_per_second_pps),                                                  //  output,   width = 1,                  master_tod_top_0_pulse_per_second.pps
		.mtod_subsys_master_tod_top_0_i_upstr_pll_lock           (mtod_subsys_master_tod_top_0_i_upstr_pll_lock),                                          //   input,   width = 1,           mtod_subsys_master_tod_top_0_i_upstr_pll.lock
		.mtod_subsys_clk100_in_clk_clk                           (sys_manager_clk_100_out_clk_clk),                                                        //   input,   width = 1,                          mtod_subsys_clk100_in_clk.clk
		.mtod_subsys_pps_load_tod_0_period_clock_clk             (sys_manager_qsys_top_master_todclk_0_out_clk_clk),                                       //   input,   width = 1,            mtod_subsys_pps_load_tod_0_period_clock.clk
		.mtod_subsys_pps_load_tod_0_reset_reset                  (rst_controller_005_reset_out_reset),                                                     //   input,   width = 1,                   mtod_subsys_pps_load_tod_0_reset.reset
		.mtod_subsys_pps_load_tod_0_csr_reset_reset              (rst_controller_005_reset_out_reset),                                                     //   input,   width = 1,               mtod_subsys_pps_load_tod_0_csr_reset.reset
		.mtod_subsys_pps_load_tod_0_csr_readdata                 (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_readdata),                 //  output,  width = 32,                     mtod_subsys_pps_load_tod_0_csr.readdata
		.mtod_subsys_pps_load_tod_0_csr_write                    (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_write),                    //   input,   width = 1,                                                   .write
		.mtod_subsys_pps_load_tod_0_csr_read                     (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_read),                     //   input,   width = 1,                                                   .read
		.mtod_subsys_pps_load_tod_0_csr_writedata                (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_writedata),                //   input,  width = 32,                                                   .writedata
		.mtod_subsys_pps_load_tod_0_csr_waitrequest              (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_waitrequest),              //  output,   width = 1,                                                   .waitrequest
		.mtod_subsys_pps_load_tod_0_csr_address                  (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_address),                  //   input,   width = 6,                                                   .address
		.mtod_subsys_pps_in_pulse_per_second                     (mtod_subsys_pps_in_pulse_per_second),                                                    //   input,   width = 1,                                 mtod_subsys_pps_in.pulse_per_second
		.mtod_subsys_pps_load_tod_0_pps_irq_irq                  (irq_mapper_receiver11_irq),                                                              //  output,   width = 1,                 mtod_subsys_pps_load_tod_0_pps_irq.irq
		.mtod_subsys_rstn_in_reset_reset_n                       (~rst_controller_reset_out_reset),                                                        //   input,   width = 1,                          mtod_subsys_rstn_in_reset.reset_n
		.tod_slave_oran_tod_stack_tx_clk_clk                     (hssi_ss_1_o_p0_clk_tx_div_clk),                                                          //   input,   width = 1,                    tod_slave_oran_tod_stack_tx_clk.clk
		.tod_slave_oran_tod_stack_rx_clk_clk                     (hssi_ss_1_o_p0_clk_rec_div_clk_signal),                                                  //   input,   width = 1,                    tod_slave_oran_tod_stack_rx_clk.clk
		.tod_slave_oran_tod_stack_todsync_sample_clk_clk         (sys_manager_ftile_iopll_todsync_sampling_outclk0_clk),                                   //   input,   width = 1,        tod_slave_oran_tod_stack_todsync_sample_clk.clk
		.tx_oran_tod_time_of_day_96b_tdata                       (tod_subsys_0_tx_oran_tod_time_of_day_96b_tdata),                                         //  output,  width = 96,                        tx_oran_tod_time_of_day_96b.tdata
		.tx_oran_tod_time_of_day_96b_tvalid                      (tod_subsys_0_tx_oran_tod_time_of_day_96b_tvalid),                                        //  output,   width = 1,                                                   .tvalid
		.rx_oran_tod_time_of_day_96b_tdata                       (tod_subsys_0_rx_oran_tod_time_of_day_96b_tdata),                                         //  output,  width = 96,                        rx_oran_tod_time_of_day_96b.tdata
		.rx_oran_tod_time_of_day_96b_tvalid                      (tod_subsys_0_rx_oran_tod_time_of_day_96b_tvalid),                                        //  output,   width = 1,                                                   .tvalid
		.tod_slave_oran_tod_stack_tx_pll_locked_lock             (tod_slave_subsys_oran_tod_stack_tx_pll_locked_lock),                                     //   input,   width = 1,             tod_slave_oran_tod_stack_tx_pll_locked.lock
		.tod_slave_port_8_tod_stack_tx_clk_clk                   (hssi_ss_1_o_p0_clk_tx_div_clk),                                                          //   input,   width = 1,                  tod_slave_port_8_tod_stack_tx_clk.clk
		.tod_slave_port_8_tod_stack_rx_clk_clk                   (hssi_ss_1_o_p0_clk_rec_div_clk_signal),                                                  //   input,   width = 1,                  tod_slave_port_8_tod_stack_rx_clk.clk
		.tod_slave_port_8_tod_stack_todsync_sample_clk_clk       (sys_manager_ftile_iopll_todsync_sampling_outclk0_clk),                                   //   input,   width = 1,      tod_slave_port_8_tod_stack_todsync_sample_clk.clk
		.tod_slave_port_8_tod_stack_tx_tod_interface_tdata       (tod_subsys_0_tod_slave_port_8_tod_stack_tx_tod_interface_tdata),                         //  output,  width = 96,        tod_slave_port_8_tod_stack_tx_tod_interface.tdata
		.tod_slave_port_8_tod_stack_tx_tod_interface_tvalid      (tod_subsys_0_tod_slave_port_8_tod_stack_tx_tod_interface_tvalid),                        //  output,   width = 1,                                                   .tvalid
		.tod_slave_port_8_tod_stack_rx_tod_interface_tdata       (tod_subsys_0_tod_slave_port_8_tod_stack_rx_tod_interface_tdata),                         //  output,  width = 96,        tod_slave_port_8_tod_stack_rx_tod_interface.tdata
		.tod_slave_port_8_tod_stack_rx_tod_interface_tvalid      (tod_subsys_0_tod_slave_port_8_tod_stack_rx_tod_interface_tvalid),                        //  output,   width = 1,                                                   .tvalid
		.tod_slave_subsys_port_8_tod_stack_tx_pll_locked_lock    (tod_slave_subsys_port_8_tod_stack_tx_pll_locked_lock),                                   //   input,   width = 1,    tod_slave_subsys_port_8_tod_stack_tx_pll_locked.lock
		.tod_slave_tod_subsys_clk_100_in_clk_clk                 (sys_manager_clk_100_out_clk_clk),                                                        //   input,   width = 1,                tod_slave_tod_subsys_clk_100_in_clk.clk
		.tod_slave_tod_subsys_mtod_clk_in_clk_clk                (sys_manager_qsys_top_master_todclk_0_out_clk_clk),                                       //   input,   width = 1,               tod_slave_tod_subsys_mtod_clk_in_clk.clk
		.tod_slave_tod_subsys_rst_100_in_reset_reset_n           (~rst_controller_002_reset_out_reset),                                                    //   input,   width = 1,              tod_slave_tod_subsys_rst_100_in_reset.reset_n
		.tod_slave_todsync_sample_plllock_split_conduit_end_lock (sys_manager_ftile_iopll_todsync_sampling_locked_lock)                                    //   input,   width = 1, tod_slave_todsync_sample_plllock_split_conduit_end.lock
	);

	qsys_top_altera_mm_interconnect_1920_pq3wixi mm_interconnect_0 (
		.hps_sub_sys_agilex_hps_h2f_axi_master_awid                                        (hps_sub_sys_agilex_hps_h2f_axi_master_awid),                                    //   input,    width = 4,                                       hps_sub_sys_agilex_hps_h2f_axi_master.awid
		.hps_sub_sys_agilex_hps_h2f_axi_master_awaddr                                      (hps_sub_sys_agilex_hps_h2f_axi_master_awaddr),                                  //   input,   width = 32,                                                                            .awaddr
		.hps_sub_sys_agilex_hps_h2f_axi_master_awlen                                       (hps_sub_sys_agilex_hps_h2f_axi_master_awlen),                                   //   input,    width = 8,                                                                            .awlen
		.hps_sub_sys_agilex_hps_h2f_axi_master_awsize                                      (hps_sub_sys_agilex_hps_h2f_axi_master_awsize),                                  //   input,    width = 3,                                                                            .awsize
		.hps_sub_sys_agilex_hps_h2f_axi_master_awburst                                     (hps_sub_sys_agilex_hps_h2f_axi_master_awburst),                                 //   input,    width = 2,                                                                            .awburst
		.hps_sub_sys_agilex_hps_h2f_axi_master_awlock                                      (hps_sub_sys_agilex_hps_h2f_axi_master_awlock),                                  //   input,    width = 1,                                                                            .awlock
		.hps_sub_sys_agilex_hps_h2f_axi_master_awcache                                     (hps_sub_sys_agilex_hps_h2f_axi_master_awcache),                                 //   input,    width = 4,                                                                            .awcache
		.hps_sub_sys_agilex_hps_h2f_axi_master_awprot                                      (hps_sub_sys_agilex_hps_h2f_axi_master_awprot),                                  //   input,    width = 3,                                                                            .awprot
		.hps_sub_sys_agilex_hps_h2f_axi_master_awvalid                                     (hps_sub_sys_agilex_hps_h2f_axi_master_awvalid),                                 //   input,    width = 1,                                                                            .awvalid
		.hps_sub_sys_agilex_hps_h2f_axi_master_awready                                     (hps_sub_sys_agilex_hps_h2f_axi_master_awready),                                 //  output,    width = 1,                                                                            .awready
		.hps_sub_sys_agilex_hps_h2f_axi_master_wdata                                       (hps_sub_sys_agilex_hps_h2f_axi_master_wdata),                                   //   input,  width = 128,                                                                            .wdata
		.hps_sub_sys_agilex_hps_h2f_axi_master_wstrb                                       (hps_sub_sys_agilex_hps_h2f_axi_master_wstrb),                                   //   input,   width = 16,                                                                            .wstrb
		.hps_sub_sys_agilex_hps_h2f_axi_master_wlast                                       (hps_sub_sys_agilex_hps_h2f_axi_master_wlast),                                   //   input,    width = 1,                                                                            .wlast
		.hps_sub_sys_agilex_hps_h2f_axi_master_wvalid                                      (hps_sub_sys_agilex_hps_h2f_axi_master_wvalid),                                  //   input,    width = 1,                                                                            .wvalid
		.hps_sub_sys_agilex_hps_h2f_axi_master_wready                                      (hps_sub_sys_agilex_hps_h2f_axi_master_wready),                                  //  output,    width = 1,                                                                            .wready
		.hps_sub_sys_agilex_hps_h2f_axi_master_bid                                         (hps_sub_sys_agilex_hps_h2f_axi_master_bid),                                     //  output,    width = 4,                                                                            .bid
		.hps_sub_sys_agilex_hps_h2f_axi_master_bresp                                       (hps_sub_sys_agilex_hps_h2f_axi_master_bresp),                                   //  output,    width = 2,                                                                            .bresp
		.hps_sub_sys_agilex_hps_h2f_axi_master_bvalid                                      (hps_sub_sys_agilex_hps_h2f_axi_master_bvalid),                                  //  output,    width = 1,                                                                            .bvalid
		.hps_sub_sys_agilex_hps_h2f_axi_master_bready                                      (hps_sub_sys_agilex_hps_h2f_axi_master_bready),                                  //   input,    width = 1,                                                                            .bready
		.hps_sub_sys_agilex_hps_h2f_axi_master_arid                                        (hps_sub_sys_agilex_hps_h2f_axi_master_arid),                                    //   input,    width = 4,                                                                            .arid
		.hps_sub_sys_agilex_hps_h2f_axi_master_araddr                                      (hps_sub_sys_agilex_hps_h2f_axi_master_araddr),                                  //   input,   width = 32,                                                                            .araddr
		.hps_sub_sys_agilex_hps_h2f_axi_master_arlen                                       (hps_sub_sys_agilex_hps_h2f_axi_master_arlen),                                   //   input,    width = 8,                                                                            .arlen
		.hps_sub_sys_agilex_hps_h2f_axi_master_arsize                                      (hps_sub_sys_agilex_hps_h2f_axi_master_arsize),                                  //   input,    width = 3,                                                                            .arsize
		.hps_sub_sys_agilex_hps_h2f_axi_master_arburst                                     (hps_sub_sys_agilex_hps_h2f_axi_master_arburst),                                 //   input,    width = 2,                                                                            .arburst
		.hps_sub_sys_agilex_hps_h2f_axi_master_arlock                                      (hps_sub_sys_agilex_hps_h2f_axi_master_arlock),                                  //   input,    width = 1,                                                                            .arlock
		.hps_sub_sys_agilex_hps_h2f_axi_master_arcache                                     (hps_sub_sys_agilex_hps_h2f_axi_master_arcache),                                 //   input,    width = 4,                                                                            .arcache
		.hps_sub_sys_agilex_hps_h2f_axi_master_arprot                                      (hps_sub_sys_agilex_hps_h2f_axi_master_arprot),                                  //   input,    width = 3,                                                                            .arprot
		.hps_sub_sys_agilex_hps_h2f_axi_master_arvalid                                     (hps_sub_sys_agilex_hps_h2f_axi_master_arvalid),                                 //   input,    width = 1,                                                                            .arvalid
		.hps_sub_sys_agilex_hps_h2f_axi_master_arready                                     (hps_sub_sys_agilex_hps_h2f_axi_master_arready),                                 //  output,    width = 1,                                                                            .arready
		.hps_sub_sys_agilex_hps_h2f_axi_master_rid                                         (hps_sub_sys_agilex_hps_h2f_axi_master_rid),                                     //  output,    width = 4,                                                                            .rid
		.hps_sub_sys_agilex_hps_h2f_axi_master_rdata                                       (hps_sub_sys_agilex_hps_h2f_axi_master_rdata),                                   //  output,  width = 128,                                                                            .rdata
		.hps_sub_sys_agilex_hps_h2f_axi_master_rresp                                       (hps_sub_sys_agilex_hps_h2f_axi_master_rresp),                                   //  output,    width = 2,                                                                            .rresp
		.hps_sub_sys_agilex_hps_h2f_axi_master_rlast                                       (hps_sub_sys_agilex_hps_h2f_axi_master_rlast),                                   //  output,    width = 1,                                                                            .rlast
		.hps_sub_sys_agilex_hps_h2f_axi_master_rvalid                                      (hps_sub_sys_agilex_hps_h2f_axi_master_rvalid),                                  //  output,    width = 1,                                                                            .rvalid
		.hps_sub_sys_agilex_hps_h2f_axi_master_rready                                      (hps_sub_sys_agilex_hps_h2f_axi_master_rready),                                  //   input,    width = 1,                                                                            .rready
		.jtg_mst_fpga_m2ocm_pb_m0_address                                                  (jtg_mst_fpga_m2ocm_pb_m0_address),                                              //   input,   width = 18,                                                    jtg_mst_fpga_m2ocm_pb_m0.address
		.jtg_mst_fpga_m2ocm_pb_m0_waitrequest                                              (jtg_mst_fpga_m2ocm_pb_m0_waitrequest),                                          //  output,    width = 1,                                                                            .waitrequest
		.jtg_mst_fpga_m2ocm_pb_m0_burstcount                                               (jtg_mst_fpga_m2ocm_pb_m0_burstcount),                                           //   input,    width = 1,                                                                            .burstcount
		.jtg_mst_fpga_m2ocm_pb_m0_byteenable                                               (jtg_mst_fpga_m2ocm_pb_m0_byteenable),                                           //   input,   width = 16,                                                                            .byteenable
		.jtg_mst_fpga_m2ocm_pb_m0_read                                                     (jtg_mst_fpga_m2ocm_pb_m0_read),                                                 //   input,    width = 1,                                                                            .read
		.jtg_mst_fpga_m2ocm_pb_m0_readdata                                                 (jtg_mst_fpga_m2ocm_pb_m0_readdata),                                             //  output,  width = 128,                                                                            .readdata
		.jtg_mst_fpga_m2ocm_pb_m0_readdatavalid                                            (jtg_mst_fpga_m2ocm_pb_m0_readdatavalid),                                        //  output,    width = 1,                                                                            .readdatavalid
		.jtg_mst_fpga_m2ocm_pb_m0_write                                                    (jtg_mst_fpga_m2ocm_pb_m0_write),                                                //   input,    width = 1,                                                                            .write
		.jtg_mst_fpga_m2ocm_pb_m0_writedata                                                (jtg_mst_fpga_m2ocm_pb_m0_writedata),                                            //   input,  width = 128,                                                                            .writedata
		.jtg_mst_fpga_m2ocm_pb_m0_debugaccess                                              (jtg_mst_fpga_m2ocm_pb_m0_debugaccess),                                          //   input,    width = 1,                                                                            .debugaccess
		.dma_subsys_dma_subsys_port8_csr_address                                           (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_address),                     //  output,    width = 8,                                             dma_subsys_dma_subsys_port8_csr.address
		.dma_subsys_dma_subsys_port8_csr_write                                             (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_write),                       //  output,    width = 1,                                                                            .write
		.dma_subsys_dma_subsys_port8_csr_read                                              (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_read),                        //  output,    width = 1,                                                                            .read
		.dma_subsys_dma_subsys_port8_csr_readdata                                          (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_readdata),                    //   input,   width = 32,                                                                            .readdata
		.dma_subsys_dma_subsys_port8_csr_writedata                                         (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_writedata),                   //  output,   width = 32,                                                                            .writedata
		.dma_subsys_dma_subsys_port8_csr_burstcount                                        (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_burstcount),                  //  output,    width = 1,                                                                            .burstcount
		.dma_subsys_dma_subsys_port8_csr_byteenable                                        (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_byteenable),                  //  output,    width = 4,                                                                            .byteenable
		.dma_subsys_dma_subsys_port8_csr_readdatavalid                                     (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_readdatavalid),               //   input,    width = 1,                                                                            .readdatavalid
		.dma_subsys_dma_subsys_port8_csr_waitrequest                                       (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_waitrequest),                 //   input,    width = 1,                                                                            .waitrequest
		.dma_subsys_dma_subsys_port8_csr_debugaccess                                       (mm_interconnect_0_dma_subsys_dma_subsys_port8_csr_debugaccess),                 //  output,    width = 1,                                                                            .debugaccess
		.dfd_subsystem_ed_synth_h2f_bridge_s0_address                                      (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_address),                //  output,   width = 28,                                        dfd_subsystem_ed_synth_h2f_bridge_s0.address
		.dfd_subsystem_ed_synth_h2f_bridge_s0_write                                        (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_write),                  //  output,    width = 1,                                                                            .write
		.dfd_subsystem_ed_synth_h2f_bridge_s0_read                                         (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_read),                   //  output,    width = 1,                                                                            .read
		.dfd_subsystem_ed_synth_h2f_bridge_s0_readdata                                     (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_readdata),               //   input,  width = 512,                                                                            .readdata
		.dfd_subsystem_ed_synth_h2f_bridge_s0_writedata                                    (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_writedata),              //  output,  width = 512,                                                                            .writedata
		.dfd_subsystem_ed_synth_h2f_bridge_s0_burstcount                                   (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_burstcount),             //  output,    width = 1,                                                                            .burstcount
		.dfd_subsystem_ed_synth_h2f_bridge_s0_byteenable                                   (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_byteenable),             //  output,   width = 64,                                                                            .byteenable
		.dfd_subsystem_ed_synth_h2f_bridge_s0_readdatavalid                                (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_readdatavalid),          //   input,    width = 1,                                                                            .readdatavalid
		.dfd_subsystem_ed_synth_h2f_bridge_s0_waitrequest                                  (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_waitrequest),            //   input,    width = 1,                                                                            .waitrequest
		.dfd_subsystem_ed_synth_h2f_bridge_s0_debugaccess                                  (mm_interconnect_0_dfd_subsystem_ed_synth_h2f_bridge_s0_debugaccess),            //  output,    width = 1,                                                                            .debugaccess
		.phipps_peak_0_h2f_bridge_s0_address                                               (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_address),                         //  output,   width = 23,                                                 phipps_peak_0_h2f_bridge_s0.address
		.phipps_peak_0_h2f_bridge_s0_write                                                 (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_write),                           //  output,    width = 1,                                                                            .write
		.phipps_peak_0_h2f_bridge_s0_read                                                  (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_read),                            //  output,    width = 1,                                                                            .read
		.phipps_peak_0_h2f_bridge_s0_readdata                                              (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_readdata),                        //   input,   width = 32,                                                                            .readdata
		.phipps_peak_0_h2f_bridge_s0_writedata                                             (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_writedata),                       //  output,   width = 32,                                                                            .writedata
		.phipps_peak_0_h2f_bridge_s0_burstcount                                            (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_burstcount),                      //  output,    width = 1,                                                                            .burstcount
		.phipps_peak_0_h2f_bridge_s0_byteenable                                            (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_byteenable),                      //  output,    width = 4,                                                                            .byteenable
		.phipps_peak_0_h2f_bridge_s0_readdatavalid                                         (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_readdatavalid),                   //   input,    width = 1,                                                                            .readdatavalid
		.phipps_peak_0_h2f_bridge_s0_waitrequest                                           (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_waitrequest),                     //   input,    width = 1,                                                                            .waitrequest
		.phipps_peak_0_h2f_bridge_s0_debugaccess                                           (mm_interconnect_0_phipps_peak_0_h2f_bridge_s0_debugaccess),                     //  output,    width = 1,                                                                            .debugaccess
		.j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_address                           (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_address),     //  output,   width = 21,                             j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr.address
		.j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_write                             (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_write),       //  output,    width = 1,                                                                            .write
		.j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_read                              (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_read),        //  output,    width = 1,                                                                            .read
		.j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_readdata                          (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_readdata),    //   input,   width = 32,                                                                            .readdata
		.j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_writedata                         (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_writedata),   //  output,   width = 32,                                                                            .writedata
		.j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_byteenable                        (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_byteenable),  //  output,    width = 4,                                                                            .byteenable
		.j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_waitrequest                       (mm_interconnect_0_j204c_f_rx_tx_ip_intel_jesd204c_f_reconfig_xcvr_waitrequest), //   input,    width = 1,                                                                            .waitrequest
		.tod_subsys_0_master_tod_top_0_csr_address                                         (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_address),                   //  output,    width = 4,                                           tod_subsys_0_master_tod_top_0_csr.address
		.tod_subsys_0_master_tod_top_0_csr_write                                           (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_write),                     //  output,    width = 1,                                                                            .write
		.tod_subsys_0_master_tod_top_0_csr_read                                            (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_read),                      //  output,    width = 1,                                                                            .read
		.tod_subsys_0_master_tod_top_0_csr_readdata                                        (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_readdata),                  //   input,   width = 32,                                                                            .readdata
		.tod_subsys_0_master_tod_top_0_csr_writedata                                       (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_writedata),                 //  output,   width = 32,                                                                            .writedata
		.tod_subsys_0_master_tod_top_0_csr_waitrequest                                     (mm_interconnect_0_tod_subsys_0_master_tod_top_0_csr_waitrequest),               //   input,    width = 1,                                                                            .waitrequest
		.tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_address                               (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_address),         //  output,    width = 6,                                 tod_subsys_0_mtod_subsys_pps_load_tod_0_csr.address
		.tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_write                                 (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_write),           //  output,    width = 1,                                                                            .write
		.tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_read                                  (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_read),            //  output,    width = 1,                                                                            .read
		.tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_readdata                              (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_readdata),        //   input,   width = 32,                                                                            .readdata
		.tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_writedata                             (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_writedata),       //  output,   width = 32,                                                                            .writedata
		.tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_waitrequest                           (mm_interconnect_0_tod_subsys_0_mtod_subsys_pps_load_tod_0_csr_waitrequest),     //   input,    width = 1,                                                                            .waitrequest
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_address                                       (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_address),                 //  output,   width = 17,                                         phipps_peak_0_pwr_mtr_h2f_bridge_s0.address
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_write                                         (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_write),                   //  output,    width = 1,                                                                            .write
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_read                                          (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_read),                    //  output,    width = 1,                                                                            .read
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdata                                      (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdata),                //   input,   width = 32,                                                                            .readdata
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_writedata                                     (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_writedata),               //  output,   width = 32,                                                                            .writedata
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_burstcount                                    (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_burstcount),              //  output,    width = 1,                                                                            .burstcount
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_byteenable                                    (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_byteenable),              //  output,    width = 4,                                                                            .byteenable
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdatavalid                                 (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_readdatavalid),           //   input,    width = 1,                                                                            .readdatavalid
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_waitrequest                                   (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_waitrequest),             //   input,    width = 1,                                                                            .waitrequest
		.phipps_peak_0_pwr_mtr_h2f_bridge_s0_debugaccess                                   (mm_interconnect_0_phipps_peak_0_pwr_mtr_h2f_bridge_s0_debugaccess),             //  output,    width = 1,                                                                            .debugaccess
		.ftile_debug_status_pio_0_s1_address                                               (mm_interconnect_0_ftile_debug_status_pio_0_s1_address),                         //  output,    width = 2,                                                 ftile_debug_status_pio_0_s1.address
		.ftile_debug_status_pio_0_s1_write                                                 (mm_interconnect_0_ftile_debug_status_pio_0_s1_write),                           //  output,    width = 1,                                                                            .write
		.ftile_debug_status_pio_0_s1_readdata                                              (mm_interconnect_0_ftile_debug_status_pio_0_s1_readdata),                        //   input,   width = 32,                                                                            .readdata
		.ftile_debug_status_pio_0_s1_writedata                                             (mm_interconnect_0_ftile_debug_status_pio_0_s1_writedata),                       //  output,   width = 32,                                                                            .writedata
		.ftile_debug_status_pio_0_s1_chipselect                                            (mm_interconnect_0_ftile_debug_status_pio_0_s1_chipselect),                      //  output,    width = 1,                                                                            .chipselect
		.ocm_s1_address                                                                    (mm_interconnect_0_ocm_s1_address),                                              //  output,   width = 14,                                                                      ocm_s1.address
		.ocm_s1_write                                                                      (mm_interconnect_0_ocm_s1_write),                                                //  output,    width = 1,                                                                            .write
		.ocm_s1_readdata                                                                   (mm_interconnect_0_ocm_s1_readdata),                                             //   input,  width = 128,                                                                            .readdata
		.ocm_s1_writedata                                                                  (mm_interconnect_0_ocm_s1_writedata),                                            //  output,  width = 128,                                                                            .writedata
		.ocm_s1_byteenable                                                                 (mm_interconnect_0_ocm_s1_byteenable),                                           //  output,   width = 16,                                                                            .byteenable
		.ocm_s1_chipselect                                                                 (mm_interconnect_0_ocm_s1_chipselect),                                           //  output,    width = 1,                                                                            .chipselect
		.ocm_s1_clken                                                                      (mm_interconnect_0_ocm_s1_clken),                                                //  output,    width = 1,                                                                            .clken
		.qsfpdd_status_pio_s1_address                                                      (mm_interconnect_0_qsfpdd_status_pio_s1_address),                                //  output,    width = 2,                                                        qsfpdd_status_pio_s1.address
		.qsfpdd_status_pio_s1_write                                                        (mm_interconnect_0_qsfpdd_status_pio_s1_write),                                  //  output,    width = 1,                                                                            .write
		.qsfpdd_status_pio_s1_readdata                                                     (mm_interconnect_0_qsfpdd_status_pio_s1_readdata),                               //   input,   width = 32,                                                                            .readdata
		.qsfpdd_status_pio_s1_writedata                                                    (mm_interconnect_0_qsfpdd_status_pio_s1_writedata),                              //  output,   width = 32,                                                                            .writedata
		.qsfpdd_status_pio_s1_chipselect                                                   (mm_interconnect_0_qsfpdd_status_pio_s1_chipselect),                             //  output,    width = 1,                                                                            .chipselect
		.sys_ctrl_pio_0_s1_address                                                         (mm_interconnect_0_sys_ctrl_pio_0_s1_address),                                   //  output,    width = 2,                                                           sys_ctrl_pio_0_s1.address
		.sys_ctrl_pio_0_s1_write                                                           (mm_interconnect_0_sys_ctrl_pio_0_s1_write),                                     //  output,    width = 1,                                                                            .write
		.sys_ctrl_pio_0_s1_readdata                                                        (mm_interconnect_0_sys_ctrl_pio_0_s1_readdata),                                  //   input,   width = 32,                                                                            .readdata
		.sys_ctrl_pio_0_s1_writedata                                                       (mm_interconnect_0_sys_ctrl_pio_0_s1_writedata),                                 //  output,   width = 32,                                                                            .writedata
		.sys_ctrl_pio_0_s1_chipselect                                                      (mm_interconnect_0_sys_ctrl_pio_0_s1_chipselect),                                //  output,    width = 1,                                                                            .chipselect
		.hssi_ss_1_axi4_lite_interface_awaddr                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awaddr),                        //  output,   width = 26,                                               hssi_ss_1_axi4_lite_interface.awaddr
		.hssi_ss_1_axi4_lite_interface_awprot                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awprot),                        //  output,    width = 3,                                                                            .awprot
		.hssi_ss_1_axi4_lite_interface_awvalid                                             (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awvalid),                       //  output,    width = 1,                                                                            .awvalid
		.hssi_ss_1_axi4_lite_interface_awready                                             (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_awready),                       //   input,    width = 1,                                                                            .awready
		.hssi_ss_1_axi4_lite_interface_wdata                                               (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wdata),                         //  output,   width = 32,                                                                            .wdata
		.hssi_ss_1_axi4_lite_interface_wstrb                                               (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wstrb),                         //  output,    width = 4,                                                                            .wstrb
		.hssi_ss_1_axi4_lite_interface_wvalid                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wvalid),                        //  output,    width = 1,                                                                            .wvalid
		.hssi_ss_1_axi4_lite_interface_wready                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_wready),                        //   input,    width = 1,                                                                            .wready
		.hssi_ss_1_axi4_lite_interface_bresp                                               (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bresp),                         //   input,    width = 2,                                                                            .bresp
		.hssi_ss_1_axi4_lite_interface_bvalid                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bvalid),                        //   input,    width = 1,                                                                            .bvalid
		.hssi_ss_1_axi4_lite_interface_bready                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_bready),                        //  output,    width = 1,                                                                            .bready
		.hssi_ss_1_axi4_lite_interface_araddr                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_araddr),                        //  output,   width = 26,                                                                            .araddr
		.hssi_ss_1_axi4_lite_interface_arprot                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arprot),                        //  output,    width = 3,                                                                            .arprot
		.hssi_ss_1_axi4_lite_interface_arvalid                                             (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arvalid),                       //  output,    width = 1,                                                                            .arvalid
		.hssi_ss_1_axi4_lite_interface_arready                                             (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_arready),                       //   input,    width = 1,                                                                            .arready
		.hssi_ss_1_axi4_lite_interface_rdata                                               (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rdata),                         //   input,   width = 32,                                                                            .rdata
		.hssi_ss_1_axi4_lite_interface_rresp                                               (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rresp),                         //   input,    width = 2,                                                                            .rresp
		.hssi_ss_1_axi4_lite_interface_rvalid                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rvalid),                        //   input,    width = 1,                                                                            .rvalid
		.hssi_ss_1_axi4_lite_interface_rready                                              (mm_interconnect_0_hssi_ss_1_axi4_lite_interface_rready),                        //  output,    width = 1,                                                                            .rready
		.hps_sub_sys_agilex_hps_h2f_axi_reset_reset_bridge_in_reset_reset                  (rst_controller_002_reset_out_reset),                                            //   input,    width = 1,                  hps_sub_sys_agilex_hps_h2f_axi_reset_reset_bridge_in_reset.reset
		.jtg_mst_reset_reset_bridge_in_reset_reset                                         (rst_controller_002_reset_out_reset),                                            //   input,    width = 1,                                         jtg_mst_reset_reset_bridge_in_reset.reset
		.dfd_subsystem_reset_csr_reset_bridge_in_reset_reset                               (rst_controller_006_reset_out_reset),                                            //   input,    width = 1,                               dfd_subsystem_reset_csr_reset_bridge_in_reset.reset
		.dfd_subsystem_ed_synth_h2f_bridge_s0_translator_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                                            //   input,    width = 1, dfd_subsystem_ed_synth_h2f_bridge_s0_translator_reset_reset_bridge_in_reset.reset
		.sys_manager_clk_100_out_clk_clk                                                   (sys_manager_clk_100_out_clk_clk),                                               //   input,    width = 1,                                                 sys_manager_clk_100_out_clk.clk
		.clk_ss_0_clk_csr_out_clk_clk                                                      (clk_ss_0_clk_csr_out_clk_clk)                                                   //   input,    width = 1,                                                    clk_ss_0_clk_csr_out_clk.clk
	);

	qsys_top_altera_mm_interconnect_1920_b6r35vi mm_interconnect_1 (
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awid                               (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awid),                                          //   input,    width = 4,                              hps_sub_sys_agilex_hps_h2f_lw_axi_master.awid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awaddr                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awaddr),                                        //   input,   width = 21,                                                                      .awaddr
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlen                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlen),                                         //   input,    width = 8,                                                                      .awlen
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awsize                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awsize),                                        //   input,    width = 3,                                                                      .awsize
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awburst                            (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awburst),                                       //   input,    width = 2,                                                                      .awburst
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlock                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awlock),                                        //   input,    width = 1,                                                                      .awlock
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awcache                            (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awcache),                                       //   input,    width = 4,                                                                      .awcache
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awprot                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awprot),                                        //   input,    width = 3,                                                                      .awprot
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awvalid                            (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awvalid),                                       //   input,    width = 1,                                                                      .awvalid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_awready                            (hps_sub_sys_agilex_hps_h2f_lw_axi_master_awready),                                       //  output,    width = 1,                                                                      .awready
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_wdata                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wdata),                                         //   input,   width = 32,                                                                      .wdata
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_wstrb                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wstrb),                                         //   input,    width = 4,                                                                      .wstrb
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_wlast                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wlast),                                         //   input,    width = 1,                                                                      .wlast
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_wvalid                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wvalid),                                        //   input,    width = 1,                                                                      .wvalid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_wready                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_wready),                                        //  output,    width = 1,                                                                      .wready
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_bid                                (hps_sub_sys_agilex_hps_h2f_lw_axi_master_bid),                                           //  output,    width = 4,                                                                      .bid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_bresp                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_bresp),                                         //  output,    width = 2,                                                                      .bresp
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_bvalid                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_bvalid),                                        //  output,    width = 1,                                                                      .bvalid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_bready                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_bready),                                        //   input,    width = 1,                                                                      .bready
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arid                               (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arid),                                          //   input,    width = 4,                                                                      .arid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_araddr                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_araddr),                                        //   input,   width = 21,                                                                      .araddr
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlen                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlen),                                         //   input,    width = 8,                                                                      .arlen
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arsize                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arsize),                                        //   input,    width = 3,                                                                      .arsize
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arburst                            (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arburst),                                       //   input,    width = 2,                                                                      .arburst
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlock                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arlock),                                        //   input,    width = 1,                                                                      .arlock
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arcache                            (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arcache),                                       //   input,    width = 4,                                                                      .arcache
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arprot                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arprot),                                        //   input,    width = 3,                                                                      .arprot
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arvalid                            (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arvalid),                                       //   input,    width = 1,                                                                      .arvalid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_arready                            (hps_sub_sys_agilex_hps_h2f_lw_axi_master_arready),                                       //  output,    width = 1,                                                                      .arready
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_rid                                (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rid),                                           //  output,    width = 4,                                                                      .rid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_rdata                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rdata),                                         //  output,   width = 32,                                                                      .rdata
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_rresp                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rresp),                                         //  output,    width = 2,                                                                      .rresp
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_rlast                              (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rlast),                                         //  output,    width = 1,                                                                      .rlast
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_rvalid                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rvalid),                                        //  output,    width = 1,                                                                      .rvalid
		.hps_sub_sys_agilex_hps_h2f_lw_axi_master_rready                             (hps_sub_sys_agilex_hps_h2f_lw_axi_master_rready),                                        //   input,    width = 1,                                                                      .rready
		.jtg_mst_fpga_m_master_address                                               (jtg_mst_fpga_m_master_address),                                                          //   input,   width = 32,                                                 jtg_mst_fpga_m_master.address
		.jtg_mst_fpga_m_master_waitrequest                                           (jtg_mst_fpga_m_master_waitrequest),                                                      //  output,    width = 1,                                                                      .waitrequest
		.jtg_mst_fpga_m_master_byteenable                                            (jtg_mst_fpga_m_master_byteenable),                                                       //   input,    width = 4,                                                                      .byteenable
		.jtg_mst_fpga_m_master_read                                                  (jtg_mst_fpga_m_master_read),                                                             //   input,    width = 1,                                                                      .read
		.jtg_mst_fpga_m_master_readdata                                              (jtg_mst_fpga_m_master_readdata),                                                         //  output,   width = 32,                                                                      .readdata
		.jtg_mst_fpga_m_master_readdatavalid                                         (jtg_mst_fpga_m_master_readdatavalid),                                                    //  output,    width = 1,                                                                      .readdatavalid
		.jtg_mst_fpga_m_master_write                                                 (jtg_mst_fpga_m_master_write),                                                            //   input,    width = 1,                                                                      .write
		.jtg_mst_fpga_m_master_writedata                                             (jtg_mst_fpga_m_master_writedata),                                                        //   input,   width = 32,                                                                      .writedata
		.hps_sub_sys_acp_0_csr_address                                               (mm_interconnect_1_hps_sub_sys_acp_0_csr_address),                                        //  output,    width = 1,                                                 hps_sub_sys_acp_0_csr.address
		.hps_sub_sys_acp_0_csr_write                                                 (mm_interconnect_1_hps_sub_sys_acp_0_csr_write),                                          //  output,    width = 1,                                                                      .write
		.hps_sub_sys_acp_0_csr_read                                                  (mm_interconnect_1_hps_sub_sys_acp_0_csr_read),                                           //  output,    width = 1,                                                                      .read
		.hps_sub_sys_acp_0_csr_readdata                                              (mm_interconnect_1_hps_sub_sys_acp_0_csr_readdata),                                       //   input,   width = 32,                                                                      .readdata
		.hps_sub_sys_acp_0_csr_writedata                                             (mm_interconnect_1_hps_sub_sys_acp_0_csr_writedata),                                      //  output,   width = 32,                                                                      .writedata
		.phipps_peak_0_h2f_lw_bridge_s0_address                                      (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_address),                               //  output,   width = 20,                                        phipps_peak_0_h2f_lw_bridge_s0.address
		.phipps_peak_0_h2f_lw_bridge_s0_write                                        (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_write),                                 //  output,    width = 1,                                                                      .write
		.phipps_peak_0_h2f_lw_bridge_s0_read                                         (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_read),                                  //  output,    width = 1,                                                                      .read
		.phipps_peak_0_h2f_lw_bridge_s0_readdata                                     (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_readdata),                              //   input,   width = 32,                                                                      .readdata
		.phipps_peak_0_h2f_lw_bridge_s0_writedata                                    (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_writedata),                             //  output,   width = 32,                                                                      .writedata
		.phipps_peak_0_h2f_lw_bridge_s0_burstcount                                   (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_burstcount),                            //  output,    width = 1,                                                                      .burstcount
		.phipps_peak_0_h2f_lw_bridge_s0_byteenable                                   (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_byteenable),                            //  output,    width = 4,                                                                      .byteenable
		.phipps_peak_0_h2f_lw_bridge_s0_readdatavalid                                (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_readdatavalid),                         //   input,    width = 1,                                                                      .readdatavalid
		.phipps_peak_0_h2f_lw_bridge_s0_waitrequest                                  (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_waitrequest),                           //   input,    width = 1,                                                                      .waitrequest
		.phipps_peak_0_h2f_lw_bridge_s0_debugaccess                                  (mm_interconnect_1_phipps_peak_0_h2f_lw_bridge_s0_debugaccess),                           //  output,    width = 1,                                                                      .debugaccess
		.dfd_subsystem_h2f_lw_bridge_s0_address                                      (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_address),                               //  output,   width = 13,                                        dfd_subsystem_h2f_lw_bridge_s0.address
		.dfd_subsystem_h2f_lw_bridge_s0_write                                        (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_write),                                 //  output,    width = 1,                                                                      .write
		.dfd_subsystem_h2f_lw_bridge_s0_read                                         (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_read),                                  //  output,    width = 1,                                                                      .read
		.dfd_subsystem_h2f_lw_bridge_s0_readdata                                     (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_readdata),                              //   input,   width = 32,                                                                      .readdata
		.dfd_subsystem_h2f_lw_bridge_s0_writedata                                    (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_writedata),                             //  output,   width = 32,                                                                      .writedata
		.dfd_subsystem_h2f_lw_bridge_s0_burstcount                                   (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_burstcount),                            //  output,    width = 1,                                                                      .burstcount
		.dfd_subsystem_h2f_lw_bridge_s0_byteenable                                   (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_byteenable),                            //  output,    width = 4,                                                                      .byteenable
		.dfd_subsystem_h2f_lw_bridge_s0_readdatavalid                                (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_readdatavalid),                         //   input,    width = 1,                                                                      .readdatavalid
		.dfd_subsystem_h2f_lw_bridge_s0_waitrequest                                  (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_waitrequest),                           //   input,    width = 1,                                                                      .waitrequest
		.dfd_subsystem_h2f_lw_bridge_s0_debugaccess                                  (mm_interconnect_1_dfd_subsystem_h2f_lw_bridge_s0_debugaccess),                           //  output,    width = 1,                                                                      .debugaccess
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_address                      (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_address),               //  output,   width = 10,                        j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs.address
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_write                        (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_write),                 //  output,    width = 1,                                                                      .write
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_read                         (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_read),                  //  output,    width = 1,                                                                      .read
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_readdata                     (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_readdata),              //   input,   width = 32,                                                                      .readdata
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_writedata                    (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_writedata),             //  output,   width = 32,                                                                      .writedata
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_waitrequest                  (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_waitrequest),           //   input,    width = 1,                                                                      .waitrequest
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_chipselect                   (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_rx_avs_chipselect),            //  output,    width = 1,                                                                      .chipselect
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_address                      (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_address),               //  output,   width = 10,                        j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs.address
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_write                        (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_write),                 //  output,    width = 1,                                                                      .write
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_read                         (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_read),                  //  output,    width = 1,                                                                      .read
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_readdata                     (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_readdata),              //   input,   width = 32,                                                                      .readdata
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_writedata                    (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_writedata),             //  output,   width = 32,                                                                      .writedata
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_waitrequest                  (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_waitrequest),           //   input,    width = 1,                                                                      .waitrequest
		.j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_chipselect                   (mm_interconnect_1_j204c_f_rx_tx_ip_intel_jesd204c_f_j204c_tx_avs_chipselect),            //  output,    width = 1,                                                                      .chipselect
		.periph_pb_cpu_0_s0_address                                                  (mm_interconnect_1_periph_pb_cpu_0_s0_address),                                           //  output,    width = 9,                                                    periph_pb_cpu_0_s0.address
		.periph_pb_cpu_0_s0_write                                                    (mm_interconnect_1_periph_pb_cpu_0_s0_write),                                             //  output,    width = 1,                                                                      .write
		.periph_pb_cpu_0_s0_read                                                     (mm_interconnect_1_periph_pb_cpu_0_s0_read),                                              //  output,    width = 1,                                                                      .read
		.periph_pb_cpu_0_s0_readdata                                                 (mm_interconnect_1_periph_pb_cpu_0_s0_readdata),                                          //   input,   width = 32,                                                                      .readdata
		.periph_pb_cpu_0_s0_writedata                                                (mm_interconnect_1_periph_pb_cpu_0_s0_writedata),                                         //  output,   width = 32,                                                                      .writedata
		.periph_pb_cpu_0_s0_burstcount                                               (mm_interconnect_1_periph_pb_cpu_0_s0_burstcount),                                        //  output,    width = 1,                                                                      .burstcount
		.periph_pb_cpu_0_s0_byteenable                                               (mm_interconnect_1_periph_pb_cpu_0_s0_byteenable),                                        //  output,    width = 4,                                                                      .byteenable
		.periph_pb_cpu_0_s0_readdatavalid                                            (mm_interconnect_1_periph_pb_cpu_0_s0_readdatavalid),                                     //   input,    width = 1,                                                                      .readdatavalid
		.periph_pb_cpu_0_s0_waitrequest                                              (mm_interconnect_1_periph_pb_cpu_0_s0_waitrequest),                                       //   input,    width = 1,                                                                      .waitrequest
		.periph_pb_cpu_0_s0_debugaccess                                              (mm_interconnect_1_periph_pb_cpu_0_s0_debugaccess),                                       //  output,    width = 1,                                                                      .debugaccess
		.j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_address                           (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_address),                    //  output,    width = 8,                             j204c_f_rx_tx_ip_reset_sequencer_0_av_csr.address
		.j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_write                             (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_write),                      //  output,    width = 1,                                                                      .write
		.j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_read                              (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_read),                       //  output,    width = 1,                                                                      .read
		.j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_readdata                          (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_readdata),                   //   input,   width = 32,                                                                      .readdata
		.j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_writedata                         (mm_interconnect_1_j204c_f_rx_tx_ip_reset_sequencer_0_av_csr_writedata),                  //  output,   width = 32,                                                                      .writedata
		.sys_manager_sysid_control_slave_address                                     (mm_interconnect_1_sys_manager_sysid_control_slave_address),                              //  output,    width = 1,                                       sys_manager_sysid_control_slave.address
		.sys_manager_sysid_control_slave_readdata                                    (mm_interconnect_1_sys_manager_sysid_control_slave_readdata),                             //   input,   width = 32,                                                                      .readdata
		.tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_address              (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_address),       //  output,    width = 5,                tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr.address
		.tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_write                (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_write),         //  output,    width = 1,                                                                      .write
		.tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_read                 (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_read),          //  output,    width = 1,                                                                      .read
		.tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata             (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata),      //   input,   width = 32,                                                                      .readdata
		.tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata            (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata),     //  output,   width = 32,                                                                      .writedata
		.tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid        (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid), //   input,    width = 1,                                                                      .readdatavalid
		.tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest          (mm_interconnect_1_tod_subsys_0_tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest),   //   input,    width = 1,                                                                      .waitrequest
		.jtg_mst_fpga_m2ocm_pb_s0_address                                            (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_address),                                     //  output,   width = 18,                                              jtg_mst_fpga_m2ocm_pb_s0.address
		.jtg_mst_fpga_m2ocm_pb_s0_write                                              (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_write),                                       //  output,    width = 1,                                                                      .write
		.jtg_mst_fpga_m2ocm_pb_s0_read                                               (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_read),                                        //  output,    width = 1,                                                                      .read
		.jtg_mst_fpga_m2ocm_pb_s0_readdata                                           (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_readdata),                                    //   input,  width = 128,                                                                      .readdata
		.jtg_mst_fpga_m2ocm_pb_s0_writedata                                          (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_writedata),                                   //  output,  width = 128,                                                                      .writedata
		.jtg_mst_fpga_m2ocm_pb_s0_burstcount                                         (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_burstcount),                                  //  output,    width = 1,                                                                      .burstcount
		.jtg_mst_fpga_m2ocm_pb_s0_byteenable                                         (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_byteenable),                                  //  output,   width = 16,                                                                      .byteenable
		.jtg_mst_fpga_m2ocm_pb_s0_readdatavalid                                      (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_readdatavalid),                               //   input,    width = 1,                                                                      .readdatavalid
		.jtg_mst_fpga_m2ocm_pb_s0_waitrequest                                        (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_waitrequest),                                 //   input,    width = 1,                                                                      .waitrequest
		.jtg_mst_fpga_m2ocm_pb_s0_debugaccess                                        (mm_interconnect_1_jtg_mst_fpga_m2ocm_pb_s0_debugaccess),                                 //  output,    width = 1,                                                                      .debugaccess
		.hps_sub_sys_agilex_hps_h2f_lw_axi_reset_reset_bridge_in_reset_reset         (rst_controller_002_reset_out_reset),                                                     //   input,    width = 1,         hps_sub_sys_agilex_hps_h2f_lw_axi_reset_reset_bridge_in_reset.reset
		.jtg_mst_reset_reset_bridge_in_reset_reset                                   (rst_controller_002_reset_out_reset),                                                     //   input,    width = 1,                                   jtg_mst_reset_reset_bridge_in_reset.reset
		.phipps_peak_0_csr_in_reset_reset_bridge_in_reset_reset                      (rst_controller_006_reset_out_reset),                                                     //   input,    width = 1,                      phipps_peak_0_csr_in_reset_reset_bridge_in_reset.reset
		.phipps_peak_0_h2f_lw_bridge_s0_translator_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                                                     //   input,    width = 1, phipps_peak_0_h2f_lw_bridge_s0_translator_reset_reset_bridge_in_reset.reset
		.sys_manager_clk_100_out_clk_clk                                             (sys_manager_clk_100_out_clk_clk),                                                        //   input,    width = 1,                                           sys_manager_clk_100_out_clk.clk
		.clk_ss_0_clk_csr_out_clk_clk                                                (clk_ss_0_clk_csr_out_clk_clk)                                                            //   input,    width = 1,                                              clk_ss_0_clk_csr_out_clk.clk
	);

	qsys_top_altera_mm_interconnect_1920_tzxrmbi mm_interconnect_2 (
		.dma_subsys_dma_ss_master_m0_address                                                      (dma_subsys_dma_ss_master_m0_address),                       //   input,   width = 37,                                                        dma_subsys_dma_ss_master_m0.address
		.dma_subsys_dma_ss_master_m0_waitrequest                                                  (dma_subsys_dma_ss_master_m0_waitrequest),                   //  output,    width = 1,                                                                                   .waitrequest
		.dma_subsys_dma_ss_master_m0_burstcount                                                   (dma_subsys_dma_ss_master_m0_burstcount),                    //   input,    width = 5,                                                                                   .burstcount
		.dma_subsys_dma_ss_master_m0_byteenable                                                   (dma_subsys_dma_ss_master_m0_byteenable),                    //   input,   width = 64,                                                                                   .byteenable
		.dma_subsys_dma_ss_master_m0_read                                                         (dma_subsys_dma_ss_master_m0_read),                          //   input,    width = 1,                                                                                   .read
		.dma_subsys_dma_ss_master_m0_readdata                                                     (dma_subsys_dma_ss_master_m0_readdata),                      //  output,  width = 512,                                                                                   .readdata
		.dma_subsys_dma_ss_master_m0_readdatavalid                                                (dma_subsys_dma_ss_master_m0_readdatavalid),                 //  output,    width = 1,                                                                                   .readdatavalid
		.dma_subsys_dma_ss_master_m0_write                                                        (dma_subsys_dma_ss_master_m0_write),                         //   input,    width = 1,                                                                                   .write
		.dma_subsys_dma_ss_master_m0_writedata                                                    (dma_subsys_dma_ss_master_m0_writedata),                     //   input,  width = 512,                                                                                   .writedata
		.dma_subsys_dma_ss_master_m0_debugaccess                                                  (dma_subsys_dma_ss_master_m0_debugaccess),                   //   input,    width = 1,                                                                                   .debugaccess
		.dma_subsys_dma_ss_master_m0_response                                                     (dma_subsys_dma_ss_master_m0_response),                      //  output,    width = 2,                                                                                   .response
		.dma_subsys_dma_ss_master_m0_writeresponsevalid                                           (dma_subsys_dma_ss_master_m0_writeresponsevalid),            //  output,    width = 1,                                                                                   .writeresponsevalid
		.dma_subsys_ext_hps_m_master_expanded_master_address                                      (dma_subsys_ext_hps_m_master_expanded_master_address),       //   input,   width = 37,                                        dma_subsys_ext_hps_m_master_expanded_master.address
		.dma_subsys_ext_hps_m_master_expanded_master_waitrequest                                  (dma_subsys_ext_hps_m_master_expanded_master_waitrequest),   //  output,    width = 1,                                                                                   .waitrequest
		.dma_subsys_ext_hps_m_master_expanded_master_burstcount                                   (dma_subsys_ext_hps_m_master_expanded_master_burstcount),    //   input,    width = 1,                                                                                   .burstcount
		.dma_subsys_ext_hps_m_master_expanded_master_byteenable                                   (dma_subsys_ext_hps_m_master_expanded_master_byteenable),    //   input,    width = 4,                                                                                   .byteenable
		.dma_subsys_ext_hps_m_master_expanded_master_read                                         (dma_subsys_ext_hps_m_master_expanded_master_read),          //   input,    width = 1,                                                                                   .read
		.dma_subsys_ext_hps_m_master_expanded_master_readdata                                     (dma_subsys_ext_hps_m_master_expanded_master_readdata),      //  output,   width = 32,                                                                                   .readdata
		.dma_subsys_ext_hps_m_master_expanded_master_readdatavalid                                (dma_subsys_ext_hps_m_master_expanded_master_readdatavalid), //  output,    width = 1,                                                                                   .readdatavalid
		.dma_subsys_ext_hps_m_master_expanded_master_write                                        (dma_subsys_ext_hps_m_master_expanded_master_write),         //   input,    width = 1,                                                                                   .write
		.dma_subsys_ext_hps_m_master_expanded_master_writedata                                    (dma_subsys_ext_hps_m_master_expanded_master_writedata),     //   input,   width = 32,                                                                                   .writedata
		.hps_sub_sys_acp_0_s0_awid                                                                (mm_interconnect_2_hps_sub_sys_acp_0_s0_awid),               //  output,    width = 4,                                                               hps_sub_sys_acp_0_s0.awid
		.hps_sub_sys_acp_0_s0_awaddr                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_awaddr),             //  output,   width = 37,                                                                                   .awaddr
		.hps_sub_sys_acp_0_s0_awlen                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_awlen),              //  output,    width = 8,                                                                                   .awlen
		.hps_sub_sys_acp_0_s0_awsize                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_awsize),             //  output,    width = 3,                                                                                   .awsize
		.hps_sub_sys_acp_0_s0_awburst                                                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_awburst),            //  output,    width = 2,                                                                                   .awburst
		.hps_sub_sys_acp_0_s0_awlock                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_awlock),             //  output,    width = 1,                                                                                   .awlock
		.hps_sub_sys_acp_0_s0_awcache                                                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_awcache),            //  output,    width = 4,                                                                                   .awcache
		.hps_sub_sys_acp_0_s0_awprot                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_awprot),             //  output,    width = 3,                                                                                   .awprot
		.hps_sub_sys_acp_0_s0_awvalid                                                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_awvalid),            //  output,    width = 1,                                                                                   .awvalid
		.hps_sub_sys_acp_0_s0_awready                                                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_awready),            //   input,    width = 1,                                                                                   .awready
		.hps_sub_sys_acp_0_s0_wdata                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_wdata),              //  output,  width = 512,                                                                                   .wdata
		.hps_sub_sys_acp_0_s0_wstrb                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_wstrb),              //  output,   width = 64,                                                                                   .wstrb
		.hps_sub_sys_acp_0_s0_wlast                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_wlast),              //  output,    width = 1,                                                                                   .wlast
		.hps_sub_sys_acp_0_s0_wvalid                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_wvalid),             //  output,    width = 1,                                                                                   .wvalid
		.hps_sub_sys_acp_0_s0_wready                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_wready),             //   input,    width = 1,                                                                                   .wready
		.hps_sub_sys_acp_0_s0_bid                                                                 (mm_interconnect_2_hps_sub_sys_acp_0_s0_bid),                //   input,    width = 4,                                                                                   .bid
		.hps_sub_sys_acp_0_s0_bresp                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_bresp),              //   input,    width = 2,                                                                                   .bresp
		.hps_sub_sys_acp_0_s0_bvalid                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_bvalid),             //   input,    width = 1,                                                                                   .bvalid
		.hps_sub_sys_acp_0_s0_bready                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_bready),             //  output,    width = 1,                                                                                   .bready
		.hps_sub_sys_acp_0_s0_arid                                                                (mm_interconnect_2_hps_sub_sys_acp_0_s0_arid),               //  output,    width = 4,                                                                                   .arid
		.hps_sub_sys_acp_0_s0_araddr                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_araddr),             //  output,   width = 37,                                                                                   .araddr
		.hps_sub_sys_acp_0_s0_arlen                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_arlen),              //  output,    width = 8,                                                                                   .arlen
		.hps_sub_sys_acp_0_s0_arsize                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_arsize),             //  output,    width = 3,                                                                                   .arsize
		.hps_sub_sys_acp_0_s0_arburst                                                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_arburst),            //  output,    width = 2,                                                                                   .arburst
		.hps_sub_sys_acp_0_s0_arlock                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_arlock),             //  output,    width = 1,                                                                                   .arlock
		.hps_sub_sys_acp_0_s0_arcache                                                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_arcache),            //  output,    width = 4,                                                                                   .arcache
		.hps_sub_sys_acp_0_s0_arprot                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_arprot),             //  output,    width = 3,                                                                                   .arprot
		.hps_sub_sys_acp_0_s0_arvalid                                                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_arvalid),            //  output,    width = 1,                                                                                   .arvalid
		.hps_sub_sys_acp_0_s0_arready                                                             (mm_interconnect_2_hps_sub_sys_acp_0_s0_arready),            //   input,    width = 1,                                                                                   .arready
		.hps_sub_sys_acp_0_s0_rid                                                                 (mm_interconnect_2_hps_sub_sys_acp_0_s0_rid),                //   input,    width = 4,                                                                                   .rid
		.hps_sub_sys_acp_0_s0_rdata                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_rdata),              //   input,  width = 512,                                                                                   .rdata
		.hps_sub_sys_acp_0_s0_rresp                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_rresp),              //   input,    width = 2,                                                                                   .rresp
		.hps_sub_sys_acp_0_s0_rlast                                                               (mm_interconnect_2_hps_sub_sys_acp_0_s0_rlast),              //   input,    width = 1,                                                                                   .rlast
		.hps_sub_sys_acp_0_s0_rvalid                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_rvalid),             //   input,    width = 1,                                                                                   .rvalid
		.hps_sub_sys_acp_0_s0_rready                                                              (mm_interconnect_2_hps_sub_sys_acp_0_s0_rready),             //  output,    width = 1,                                                                                   .rready
		.dma_subsys_dma_rst_100_in_reset_reset_bridge_in_reset_reset                              (rst_controller_007_reset_out_reset),                        //   input,    width = 1,                              dma_subsys_dma_rst_100_in_reset_reset_bridge_in_reset.reset
		.hps_sub_sys_acp_0_reset_reset_bridge_in_reset_reset                                      (rst_controller_008_reset_out_reset),                        //   input,    width = 1,                                      hps_sub_sys_acp_0_reset_reset_bridge_in_reset.reset
		.dma_subsys_dma_ss_master_m0_translator_reset_reset_bridge_in_reset_reset                 (rst_controller_007_reset_out_reset),                        //   input,    width = 1,                 dma_subsys_dma_ss_master_m0_translator_reset_reset_bridge_in_reset.reset
		.dma_subsys_ext_hps_m_master_expanded_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                        //   input,    width = 1, dma_subsys_ext_hps_m_master_expanded_master_translator_reset_reset_bridge_in_reset.reset
		.hps_sub_sys_acp_0_s0_translator_clk_reset_reset_bridge_in_reset_reset                    (rst_controller_008_reset_out_reset),                        //   input,    width = 1,                    hps_sub_sys_acp_0_s0_translator_clk_reset_reset_bridge_in_reset.reset
		.crosser_002_in_clk_reset_reset_bridge_in_reset_reset                                     (rst_controller_002_reset_out_reset),                        //   input,    width = 1,                                     crosser_002_in_clk_reset_reset_bridge_in_reset.reset
		.dma_subsys_dma_clk_out_bridge_0_out_clk_clk                                              (dma_subsys_dma_clk_out_bridge_0_out_clk_clk),               //   input,    width = 1,                                            dma_subsys_dma_clk_out_bridge_0_out_clk.clk
		.sys_manager_clk_100_out_clk_clk                                                          (sys_manager_clk_100_out_clk_clk),                           //   input,    width = 1,                                                        sys_manager_clk_100_out_clk.clk
		.dma_subsys_acp_bridge_in_clk_clk                                                         (dma_subsys_acp_bridge_in_clk_clk)                           //   input,    width = 1,                                                       dma_subsys_acp_bridge_in_clk.clk
	);

	qsys_top_altera_mm_interconnect_1920_j7dvj2y mm_interconnect_3 (
		.jtg_mst_hps_m_master_address                             (jtg_mst_hps_m_master_address),                                               //   input,  width = 32,                       jtg_mst_hps_m_master.address
		.jtg_mst_hps_m_master_waitrequest                         (jtg_mst_hps_m_master_waitrequest),                                           //  output,   width = 1,                                           .waitrequest
		.jtg_mst_hps_m_master_byteenable                          (jtg_mst_hps_m_master_byteenable),                                            //   input,   width = 4,                                           .byteenable
		.jtg_mst_hps_m_master_read                                (jtg_mst_hps_m_master_read),                                                  //   input,   width = 1,                                           .read
		.jtg_mst_hps_m_master_readdata                            (jtg_mst_hps_m_master_readdata),                                              //  output,  width = 32,                                           .readdata
		.jtg_mst_hps_m_master_readdatavalid                       (jtg_mst_hps_m_master_readdatavalid),                                         //  output,   width = 1,                                           .readdatavalid
		.jtg_mst_hps_m_master_write                               (jtg_mst_hps_m_master_write),                                                 //   input,   width = 1,                                           .write
		.jtg_mst_hps_m_master_writedata                           (jtg_mst_hps_m_master_writedata),                                             //   input,  width = 32,                                           .writedata
		.dma_subsys_ext_hps_m_master_windowed_slave_address       (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_address),       //  output,  width = 30, dma_subsys_ext_hps_m_master_windowed_slave.address
		.dma_subsys_ext_hps_m_master_windowed_slave_write         (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_write),         //  output,   width = 1,                                           .write
		.dma_subsys_ext_hps_m_master_windowed_slave_read          (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_read),          //  output,   width = 1,                                           .read
		.dma_subsys_ext_hps_m_master_windowed_slave_readdata      (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_readdata),      //   input,  width = 32,                                           .readdata
		.dma_subsys_ext_hps_m_master_windowed_slave_writedata     (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_writedata),     //  output,  width = 32,                                           .writedata
		.dma_subsys_ext_hps_m_master_windowed_slave_burstcount    (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_burstcount),    //  output,   width = 1,                                           .burstcount
		.dma_subsys_ext_hps_m_master_windowed_slave_byteenable    (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_byteenable),    //  output,   width = 4,                                           .byteenable
		.dma_subsys_ext_hps_m_master_windowed_slave_readdatavalid (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_readdatavalid), //   input,   width = 1,                                           .readdatavalid
		.dma_subsys_ext_hps_m_master_windowed_slave_waitrequest   (mm_interconnect_3_dma_subsys_ext_hps_m_master_windowed_slave_waitrequest),   //   input,   width = 1,                                           .waitrequest
		.jtg_mst_reset_reset_bridge_in_reset_reset                (rst_controller_002_reset_out_reset),                                         //   input,   width = 1,        jtg_mst_reset_reset_bridge_in_reset.reset
		.sys_manager_clk_100_out_clk_clk                          (sys_manager_clk_100_out_clk_clk)                                             //   input,   width = 1,                sys_manager_clk_100_out_clk.clk
	);

	qsys_top_altera_irq_mapper_2001_rxikitq irq_mapper (
		.clk            (),                                    //   input,   width = 1,        clk.clk
		.reset          (),                                    //   input,   width = 1,  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),            //   input,   width = 1,  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),            //   input,   width = 1,  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),            //   input,   width = 1,  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),            //   input,   width = 1,  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),            //   input,   width = 1,  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),            //   input,   width = 1,  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),            //   input,   width = 1,  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),            //   input,   width = 1,  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),            //   input,   width = 1,  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),            //   input,   width = 1,  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),           //   input,   width = 1, receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq),           //   input,   width = 1, receiver11.irq
		.receiver12_irq (irq_mapper_receiver12_irq),           //   input,   width = 1, receiver12.irq
		.receiver13_irq (irq_mapper_receiver13_irq),           //   input,   width = 1, receiver13.irq
		.sender_irq     (hps_sub_sys_agilex_hps_f2h_irq0_irq)  //  output,  width = 32,     sender.irq
	);

	qsys_top_altera_irq_mapper_2001_j4mn3ji irq_mapper_001 (
		.clk           (sys_manager_clk_100_out_clk_clk), //   input,  width = 1,       clk.clk
		.reset         (rst_controller_reset_out_reset),  //   input,  width = 1, clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),        //   input,  width = 1, receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),        //   input,  width = 1, receiver1.irq
		.sender_irq    (periph_ilc_irq_irq)               //  output,  width = 2,    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~sys_manager_rst_in_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (sys_manager_clk_100_out_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_in1      (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~sys_manager_rst_in_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (dma_subsys_acp_bridge_in_clk_clk),    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                    // (terminated),                       
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_in1      (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~sys_manager_rst_in_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (sys_manager_clk_100_out_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                    // (terminated),                       
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_in1      (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~sys_manager_rst_in_out_reset_reset),   //   input,  width = 1, reset_in0.reset
		.clk            (hssi_ss_1_o_p0_clk_rec_div_clk_signal), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),    //  output,  width = 1, reset_out.reset
		.reset_req      (),                                      // (terminated),                       
		.reset_req_in0  (1'b0),                                  // (terminated),                       
		.reset_in1      (1'b0),                                  // (terminated),                       
		.reset_req_in1  (1'b0),                                  // (terminated),                       
		.reset_in2      (1'b0),                                  // (terminated),                       
		.reset_req_in2  (1'b0),                                  // (terminated),                       
		.reset_in3      (1'b0),                                  // (terminated),                       
		.reset_req_in3  (1'b0),                                  // (terminated),                       
		.reset_in4      (1'b0),                                  // (terminated),                       
		.reset_req_in4  (1'b0),                                  // (terminated),                       
		.reset_in5      (1'b0),                                  // (terminated),                       
		.reset_req_in5  (1'b0),                                  // (terminated),                       
		.reset_in6      (1'b0),                                  // (terminated),                       
		.reset_req_in6  (1'b0),                                  // (terminated),                       
		.reset_in7      (1'b0),                                  // (terminated),                       
		.reset_req_in7  (1'b0),                                  // (terminated),                       
		.reset_in8      (1'b0),                                  // (terminated),                       
		.reset_req_in8  (1'b0),                                  // (terminated),                       
		.reset_in9      (1'b0),                                  // (terminated),                       
		.reset_req_in9  (1'b0),                                  // (terminated),                       
		.reset_in10     (1'b0),                                  // (terminated),                       
		.reset_req_in10 (1'b0),                                  // (terminated),                       
		.reset_in11     (1'b0),                                  // (terminated),                       
		.reset_req_in11 (1'b0),                                  // (terminated),                       
		.reset_in12     (1'b0),                                  // (terminated),                       
		.reset_req_in12 (1'b0),                                  // (terminated),                       
		.reset_in13     (1'b0),                                  // (terminated),                       
		.reset_req_in13 (1'b0),                                  // (terminated),                       
		.reset_in14     (1'b0),                                  // (terminated),                       
		.reset_req_in14 (1'b0),                                  // (terminated),                       
		.reset_in15     (1'b0),                                  // (terminated),                       
		.reset_req_in15 (1'b0)                                   // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~sys_manager_rst_in_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (hssi_ss_1_o_p0_clk_tx_div_clk),       //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                    // (terminated),                       
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_in1      (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~sys_manager_rst_in_out_reset_reset),              //   input,  width = 1, reset_in0.reset
		.clk            (sys_manager_qsys_top_master_todclk_0_out_clk_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),               //  output,  width = 1, reset_out.reset
		.reset_req      (),                                                 // (terminated),                       
		.reset_req_in0  (1'b0),                                             // (terminated),                       
		.reset_in1      (1'b0),                                             // (terminated),                       
		.reset_req_in1  (1'b0),                                             // (terminated),                       
		.reset_in2      (1'b0),                                             // (terminated),                       
		.reset_req_in2  (1'b0),                                             // (terminated),                       
		.reset_in3      (1'b0),                                             // (terminated),                       
		.reset_req_in3  (1'b0),                                             // (terminated),                       
		.reset_in4      (1'b0),                                             // (terminated),                       
		.reset_req_in4  (1'b0),                                             // (terminated),                       
		.reset_in5      (1'b0),                                             // (terminated),                       
		.reset_req_in5  (1'b0),                                             // (terminated),                       
		.reset_in6      (1'b0),                                             // (terminated),                       
		.reset_req_in6  (1'b0),                                             // (terminated),                       
		.reset_in7      (1'b0),                                             // (terminated),                       
		.reset_req_in7  (1'b0),                                             // (terminated),                       
		.reset_in8      (1'b0),                                             // (terminated),                       
		.reset_req_in8  (1'b0),                                             // (terminated),                       
		.reset_in9      (1'b0),                                             // (terminated),                       
		.reset_req_in9  (1'b0),                                             // (terminated),                       
		.reset_in10     (1'b0),                                             // (terminated),                       
		.reset_req_in10 (1'b0),                                             // (terminated),                       
		.reset_in11     (1'b0),                                             // (terminated),                       
		.reset_req_in11 (1'b0),                                             // (terminated),                       
		.reset_in12     (1'b0),                                             // (terminated),                       
		.reset_req_in12 (1'b0),                                             // (terminated),                       
		.reset_in13     (1'b0),                                             // (terminated),                       
		.reset_req_in13 (1'b0),                                             // (terminated),                       
		.reset_in14     (1'b0),                                             // (terminated),                       
		.reset_req_in14 (1'b0),                                             // (terminated),                       
		.reset_in15     (1'b0),                                             // (terminated),                       
		.reset_req_in15 (1'b0)                                              // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~rst_ss_0_rst_csr_out_reset_reset),  //   input,  width = 1, reset_in0.reset
		.clk            (clk_ss_0_clk_csr_out_clk_clk),       //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~sys_manager_rst_in_out_reset_reset),         //   input,  width = 1, reset_in0.reset
		.clk            (dma_subsys_dma_clk_out_bridge_0_out_clk_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset),          //  output,  width = 1, reset_out.reset
		.reset_req      (),                                            // (terminated),                       
		.reset_req_in0  (1'b0),                                        // (terminated),                       
		.reset_in1      (1'b0),                                        // (terminated),                       
		.reset_req_in1  (1'b0),                                        // (terminated),                       
		.reset_in2      (1'b0),                                        // (terminated),                       
		.reset_req_in2  (1'b0),                                        // (terminated),                       
		.reset_in3      (1'b0),                                        // (terminated),                       
		.reset_req_in3  (1'b0),                                        // (terminated),                       
		.reset_in4      (1'b0),                                        // (terminated),                       
		.reset_req_in4  (1'b0),                                        // (terminated),                       
		.reset_in5      (1'b0),                                        // (terminated),                       
		.reset_req_in5  (1'b0),                                        // (terminated),                       
		.reset_in6      (1'b0),                                        // (terminated),                       
		.reset_req_in6  (1'b0),                                        // (terminated),                       
		.reset_in7      (1'b0),                                        // (terminated),                       
		.reset_req_in7  (1'b0),                                        // (terminated),                       
		.reset_in8      (1'b0),                                        // (terminated),                       
		.reset_req_in8  (1'b0),                                        // (terminated),                       
		.reset_in9      (1'b0),                                        // (terminated),                       
		.reset_req_in9  (1'b0),                                        // (terminated),                       
		.reset_in10     (1'b0),                                        // (terminated),                       
		.reset_req_in10 (1'b0),                                        // (terminated),                       
		.reset_in11     (1'b0),                                        // (terminated),                       
		.reset_req_in11 (1'b0),                                        // (terminated),                       
		.reset_in12     (1'b0),                                        // (terminated),                       
		.reset_req_in12 (1'b0),                                        // (terminated),                       
		.reset_in13     (1'b0),                                        // (terminated),                       
		.reset_req_in13 (1'b0),                                        // (terminated),                       
		.reset_in14     (1'b0),                                        // (terminated),                       
		.reset_req_in14 (1'b0),                                        // (terminated),                       
		.reset_in15     (1'b0),                                        // (terminated),                       
		.reset_req_in15 (1'b0)                                         // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~sys_manager_rst_in_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (dma_subsys_acp_bridge_in_clk_clk),    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                    // (terminated),                       
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_in1      (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

endmodule
