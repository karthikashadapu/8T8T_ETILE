// subsys_ftile_25gbe_rx_dma.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module subsys_ftile_25gbe_rx_dma (
		input  wire         dma_clk_clk,                                //                 dma_clk.clk
		output wire         csr_waitrequest,                            //                     csr.waitrequest
		output wire [31:0]  csr_readdata,                               //                        .readdata
		output wire         csr_readdatavalid,                          //                        .readdatavalid
		input  wire [0:0]   csr_burstcount,                             //                        .burstcount
		input  wire [31:0]  csr_writedata,                              //                        .writedata
		input  wire [5:0]   csr_address,                                //                        .address
		input  wire         csr_write,                                  //                        .write
		input  wire         csr_read,                                   //                        .read
		input  wire [3:0]   csr_byteenable,                             //                        .byteenable
		input  wire         csr_debugaccess,                            //                        .debugaccess
		input  wire         pktin_startofpacket,                        //                   pktin.startofpacket
		input  wire         pktin_valid,                                //                        .valid
		input  wire         pktin_endofpacket,                          //                        .endofpacket
		input  wire [63:0]  pktin_data,                                 //                        .data
		input  wire [2:0]   pktin_empty,                                //                        .empty
		input  wire [5:0]   pktin_error,                                //                        .error
		input  wire         rx_dma_fifo_0_in_ts_valid,                  //     rx_dma_fifo_0_in_ts.valid
		input  wire [95:0]  rx_dma_fifo_0_in_ts_data,                   //                        .data
		input  wire         ftile_clk_clk,                              //               ftile_clk.clk
		output wire [36:0]  prefetcher_read_master_address,             //  prefetcher_read_master.address
		output wire         prefetcher_read_master_read,                //                        .read
		input  wire [127:0] prefetcher_read_master_readdata,            //                        .readdata
		input  wire         prefetcher_read_master_waitrequest,         //                        .waitrequest
		input  wire         prefetcher_read_master_readdatavalid,       //                        .readdatavalid
		output wire [2:0]   prefetcher_read_master_burstcount,          //                        .burstcount
		output wire [36:0]  prefetcher_write_master_address,            // prefetcher_write_master.address
		output wire         prefetcher_write_master_write,              //                        .write
		output wire [15:0]  prefetcher_write_master_byteenable,         //                        .byteenable
		output wire [127:0] prefetcher_write_master_writedata,          //                        .writedata
		input  wire         prefetcher_write_master_waitrequest,        //                        .waitrequest
		input  wire [1:0]   prefetcher_write_master_response,           //                        .response
		input  wire         prefetcher_write_master_writeresponsevalid, //                        .writeresponsevalid
		output wire         irq_irq,                                    //                     irq.irq
		input  wire         reset_reset_n,                              //                   reset.reset_n
		output wire [36:0]  write_master_address,                       //            write_master.address
		output wire         write_master_write,                         //                        .write
		output wire [15:0]  write_master_byteenable,                    //                        .byteenable
		output wire [127:0] write_master_writedata,                     //                        .writedata
		input  wire         write_master_waitrequest,                   //                        .waitrequest
		output wire [4:0]   write_master_burstcount,                    //                        .burstcount
		input  wire [1:0]   write_master_response,                      //                        .response
		input  wire         write_master_writeresponsevalid             //                        .writeresponsevalid
	);

	wire          rx_dma_prefetcher_descriptor_write_dispatcher_source_valid; // rx_dma_prefetcher:st_src_descr_valid -> rx_dma_dispatcher:snk_descriptor_valid
	wire  [255:0] rx_dma_prefetcher_descriptor_write_dispatcher_source_data;  // rx_dma_prefetcher:st_src_descr_data -> rx_dma_dispatcher:snk_descriptor_data
	wire          rx_dma_prefetcher_descriptor_write_dispatcher_source_ready; // rx_dma_dispatcher:snk_descriptor_ready -> rx_dma_prefetcher:st_src_descr_ready
	wire          rx_dma_write_master_response_source_valid;                  // rx_dma_write_master:src_response_valid -> rx_dma_dispatcher:snk_write_master_valid
	wire  [255:0] rx_dma_write_master_response_source_data;                   // rx_dma_write_master:src_response_data -> rx_dma_dispatcher:snk_write_master_data
	wire          rx_dma_write_master_response_source_ready;                  // rx_dma_dispatcher:snk_write_master_ready -> rx_dma_write_master:src_response_ready
	wire          rx_dma_dispatcher_response_source_valid;                    // rx_dma_dispatcher:src_response_valid -> rx_dma_fifo_0:in_ts_resp_valid
	wire  [255:0] rx_dma_dispatcher_response_source_data;                     // rx_dma_dispatcher:src_response_data -> rx_dma_fifo_0:in_ts_resp_data
	wire          rx_dma_dispatcher_response_source_ready;                    // rx_dma_fifo_0:in_ts_resp_ready -> rx_dma_dispatcher:src_response_ready
	wire          rx_dma_dispatcher_write_command_source_valid;               // rx_dma_dispatcher:src_write_master_valid -> rx_dma_write_master:snk_command_valid
	wire  [255:0] rx_dma_dispatcher_write_command_source_data;                // rx_dma_dispatcher:src_write_master_data -> rx_dma_write_master:snk_command_data
	wire          rx_dma_dispatcher_write_command_source_ready;               // rx_dma_write_master:snk_command_ready -> rx_dma_dispatcher:src_write_master_ready
	wire          rx_dma_fifo_0_out_ts_resp_valid;                            // rx_dma_fifo_0:out_ts_resp_valid -> rx_dma_prefetcher:st_snk_valid
	wire  [255:0] rx_dma_fifo_0_out_ts_resp_data;                             // rx_dma_fifo_0:out_ts_resp_data -> rx_dma_prefetcher:st_snk_data
	wire          rx_dma_fifo_0_out_ts_resp_ready;                            // rx_dma_prefetcher:st_snk_ready -> rx_dma_fifo_0:out_ts_resp_ready
	wire          rx_dma_clock_out_clk_clk;                                   // rx_dma_clock:out_clk -> [avalon_st_adapter:in_clk_0_clk, mm_interconnect_0:rx_dma_clock_out_clk_clk, rx_dma_csr:clk, rx_dma_dispatcher:clk, rx_dma_fifo_0:csr_clk, rx_dma_fifo_0:out_st_clk, rx_dma_prefetcher:clk, rx_dma_reset:clk, rx_dma_write_master:clk]
	wire          rx_dma_ftile_clock_out_clk_clk;                             // rx_dma_ftile_clock:out_clk -> [ftile_clk_reset:clk, rst_controller:clk, rst_controller_001:clk, rx_dma_fifo_0:in_st_clk]
	wire          rx_dma_reset_out_reset_reset;                               // rx_dma_reset:out_reset_n -> [avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:rx_dma_csr_reset_reset_bridge_in_reset_reset, mm_interconnect_0:rx_dma_dispatcher_clock_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in0, rx_dma_csr:reset, rx_dma_dispatcher:reset, rx_dma_fifo_0:out_st_rst, rx_dma_prefetcher:reset, rx_dma_write_master:reset]
	wire          ftile_clk_reset_out_reset_reset;                            // ftile_clk_reset:out_reset_n -> rx_dma_fifo_0:in_st_rst
	wire          rx_dma_csr_m0_waitrequest;                                  // mm_interconnect_0:rx_dma_csr_m0_waitrequest -> rx_dma_csr:m0_waitrequest
	wire   [31:0] rx_dma_csr_m0_readdata;                                     // mm_interconnect_0:rx_dma_csr_m0_readdata -> rx_dma_csr:m0_readdata
	wire          rx_dma_csr_m0_debugaccess;                                  // rx_dma_csr:m0_debugaccess -> mm_interconnect_0:rx_dma_csr_m0_debugaccess
	wire    [5:0] rx_dma_csr_m0_address;                                      // rx_dma_csr:m0_address -> mm_interconnect_0:rx_dma_csr_m0_address
	wire          rx_dma_csr_m0_read;                                         // rx_dma_csr:m0_read -> mm_interconnect_0:rx_dma_csr_m0_read
	wire    [3:0] rx_dma_csr_m0_byteenable;                                   // rx_dma_csr:m0_byteenable -> mm_interconnect_0:rx_dma_csr_m0_byteenable
	wire          rx_dma_csr_m0_readdatavalid;                                // mm_interconnect_0:rx_dma_csr_m0_readdatavalid -> rx_dma_csr:m0_readdatavalid
	wire   [31:0] rx_dma_csr_m0_writedata;                                    // rx_dma_csr:m0_writedata -> mm_interconnect_0:rx_dma_csr_m0_writedata
	wire          rx_dma_csr_m0_write;                                        // rx_dma_csr:m0_write -> mm_interconnect_0:rx_dma_csr_m0_write
	wire    [0:0] rx_dma_csr_m0_burstcount;                                   // rx_dma_csr:m0_burstcount -> mm_interconnect_0:rx_dma_csr_m0_burstcount
	wire   [31:0] mm_interconnect_0_rx_dma_dispatcher_csr_readdata;           // rx_dma_dispatcher:csr_readdata -> mm_interconnect_0:rx_dma_dispatcher_CSR_readdata
	wire    [2:0] mm_interconnect_0_rx_dma_dispatcher_csr_address;            // mm_interconnect_0:rx_dma_dispatcher_CSR_address -> rx_dma_dispatcher:csr_address
	wire          mm_interconnect_0_rx_dma_dispatcher_csr_read;               // mm_interconnect_0:rx_dma_dispatcher_CSR_read -> rx_dma_dispatcher:csr_read
	wire    [3:0] mm_interconnect_0_rx_dma_dispatcher_csr_byteenable;         // mm_interconnect_0:rx_dma_dispatcher_CSR_byteenable -> rx_dma_dispatcher:csr_byteenable
	wire          mm_interconnect_0_rx_dma_dispatcher_csr_write;              // mm_interconnect_0:rx_dma_dispatcher_CSR_write -> rx_dma_dispatcher:csr_write
	wire   [31:0] mm_interconnect_0_rx_dma_dispatcher_csr_writedata;          // mm_interconnect_0:rx_dma_dispatcher_CSR_writedata -> rx_dma_dispatcher:csr_writedata
	wire   [31:0] mm_interconnect_0_rx_dma_prefetcher_csr_readdata;           // rx_dma_prefetcher:mm_csr_readdata -> mm_interconnect_0:rx_dma_prefetcher_Csr_readdata
	wire    [2:0] mm_interconnect_0_rx_dma_prefetcher_csr_address;            // mm_interconnect_0:rx_dma_prefetcher_Csr_address -> rx_dma_prefetcher:mm_csr_address
	wire          mm_interconnect_0_rx_dma_prefetcher_csr_read;               // mm_interconnect_0:rx_dma_prefetcher_Csr_read -> rx_dma_prefetcher:mm_csr_read
	wire          mm_interconnect_0_rx_dma_prefetcher_csr_write;              // mm_interconnect_0:rx_dma_prefetcher_Csr_write -> rx_dma_prefetcher:mm_csr_write
	wire   [31:0] mm_interconnect_0_rx_dma_prefetcher_csr_writedata;          // mm_interconnect_0:rx_dma_prefetcher_Csr_writedata -> rx_dma_prefetcher:mm_csr_writedata
	wire          rx_dma_fifo_0_out_avst_valid;                               // rx_dma_fifo_0:out_st_valid -> avalon_st_adapter:in_0_valid
	wire   [63:0] rx_dma_fifo_0_out_avst_data;                                // rx_dma_fifo_0:out_st_data -> avalon_st_adapter:in_0_data
	wire          rx_dma_fifo_0_out_avst_ready;                               // avalon_st_adapter:in_0_ready -> rx_dma_fifo_0:out_st_ready
	wire          rx_dma_fifo_0_out_avst_startofpacket;                       // rx_dma_fifo_0:out_st_sop -> avalon_st_adapter:in_0_startofpacket
	wire          rx_dma_fifo_0_out_avst_endofpacket;                         // rx_dma_fifo_0:out_st_eop -> avalon_st_adapter:in_0_endofpacket
	wire    [5:0] rx_dma_fifo_0_out_avst_error;                               // rx_dma_fifo_0:out_st_error -> avalon_st_adapter:in_0_error
	wire    [2:0] rx_dma_fifo_0_out_avst_empty;                               // rx_dma_fifo_0:out_st_empty -> avalon_st_adapter:in_0_empty
	wire          avalon_st_adapter_out_0_valid;                              // avalon_st_adapter:out_0_valid -> rx_dma_write_master:snk_valid
	wire  [127:0] avalon_st_adapter_out_0_data;                               // avalon_st_adapter:out_0_data -> rx_dma_write_master:snk_data
	wire          avalon_st_adapter_out_0_ready;                              // rx_dma_write_master:snk_ready -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                      // avalon_st_adapter:out_0_startofpacket -> rx_dma_write_master:snk_sop
	wire          avalon_st_adapter_out_0_endofpacket;                        // avalon_st_adapter:out_0_endofpacket -> rx_dma_write_master:snk_eop
	wire    [5:0] avalon_st_adapter_out_0_error;                              // avalon_st_adapter:out_0_error -> rx_dma_write_master:snk_error
	wire    [3:0] avalon_st_adapter_out_0_empty;                              // avalon_st_adapter:out_0_empty -> rx_dma_write_master:snk_empty
	wire          rst_controller_reset_out_reset;                             // rst_controller:reset_out -> ftile_clk_reset:in_reset_n
	wire          rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> rx_dma_fifo_0:csr_rst

	ftile_clk_reset ftile_clk_reset (
		.clk         (rx_dma_ftile_clock_out_clk_clk),  //   input,  width = 1,       clk.clk
		.in_reset_n  (~rst_controller_reset_out_reset), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (ftile_clk_reset_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	rx_dma_clock rx_dma_clock (
		.in_clk  (dma_clk_clk),              //   input,  width = 1,  in_clk.clk
		.out_clk (rx_dma_clock_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	rx_dma_csr rx_dma_csr (
		.clk              (rx_dma_clock_out_clk_clk),      //   input,   width = 1,   clk.clk
		.reset            (~rx_dma_reset_out_reset_reset), //   input,   width = 1, reset.reset
		.s0_waitrequest   (csr_waitrequest),               //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (csr_readdata),                  //  output,  width = 32,      .readdata
		.s0_readdatavalid (csr_readdatavalid),             //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (csr_burstcount),                //   input,   width = 1,      .burstcount
		.s0_writedata     (csr_writedata),                 //   input,  width = 32,      .writedata
		.s0_address       (csr_address),                   //   input,   width = 6,      .address
		.s0_write         (csr_write),                     //   input,   width = 1,      .write
		.s0_read          (csr_read),                      //   input,   width = 1,      .read
		.s0_byteenable    (csr_byteenable),                //   input,   width = 4,      .byteenable
		.s0_debugaccess   (csr_debugaccess),               //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (rx_dma_csr_m0_waitrequest),     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (rx_dma_csr_m0_readdata),        //   input,  width = 32,      .readdata
		.m0_readdatavalid (rx_dma_csr_m0_readdatavalid),   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (rx_dma_csr_m0_burstcount),      //  output,   width = 1,      .burstcount
		.m0_writedata     (rx_dma_csr_m0_writedata),       //  output,  width = 32,      .writedata
		.m0_address       (rx_dma_csr_m0_address),         //  output,   width = 6,      .address
		.m0_write         (rx_dma_csr_m0_write),           //  output,   width = 1,      .write
		.m0_read          (rx_dma_csr_m0_read),            //  output,   width = 1,      .read
		.m0_byteenable    (rx_dma_csr_m0_byteenable),      //  output,   width = 4,      .byteenable
		.m0_debugaccess   (rx_dma_csr_m0_debugaccess)      //  output,   width = 1,      .debugaccess
	);

	rx_dma_dispatcher rx_dma_dispatcher (
		.clk                    (rx_dma_clock_out_clk_clk),                                   //   input,    width = 1,                clock.clk
		.reset                  (~rx_dma_reset_out_reset_reset),                              //   input,    width = 1,          clock_reset.reset
		.csr_writedata          (mm_interconnect_0_rx_dma_dispatcher_csr_writedata),          //   input,   width = 32,                  CSR.writedata
		.csr_write              (mm_interconnect_0_rx_dma_dispatcher_csr_write),              //   input,    width = 1,                     .write
		.csr_byteenable         (mm_interconnect_0_rx_dma_dispatcher_csr_byteenable),         //   input,    width = 4,                     .byteenable
		.csr_readdata           (mm_interconnect_0_rx_dma_dispatcher_csr_readdata),           //  output,   width = 32,                     .readdata
		.csr_read               (mm_interconnect_0_rx_dma_dispatcher_csr_read),               //   input,    width = 1,                     .read
		.csr_address            (mm_interconnect_0_rx_dma_dispatcher_csr_address),            //   input,    width = 3,                     .address
		.src_response_data      (rx_dma_dispatcher_response_source_data),                     //  output,  width = 256,      Response_Source.data
		.src_response_valid     (rx_dma_dispatcher_response_source_valid),                    //  output,    width = 1,                     .valid
		.src_response_ready     (rx_dma_dispatcher_response_source_ready),                    //   input,    width = 1,                     .ready
		.snk_descriptor_data    (rx_dma_prefetcher_descriptor_write_dispatcher_source_data),  //   input,  width = 256,      Descriptor_Sink.data
		.snk_descriptor_valid   (rx_dma_prefetcher_descriptor_write_dispatcher_source_valid), //   input,    width = 1,                     .valid
		.snk_descriptor_ready   (rx_dma_prefetcher_descriptor_write_dispatcher_source_ready), //  output,    width = 1,                     .ready
		.src_write_master_data  (rx_dma_dispatcher_write_command_source_data),                //  output,  width = 256, Write_Command_Source.data
		.src_write_master_valid (rx_dma_dispatcher_write_command_source_valid),               //  output,    width = 1,                     .valid
		.src_write_master_ready (rx_dma_dispatcher_write_command_source_ready),               //   input,    width = 1,                     .ready
		.snk_write_master_data  (rx_dma_write_master_response_source_data),                   //   input,  width = 256,  Write_Response_Sink.data
		.snk_write_master_valid (rx_dma_write_master_response_source_valid),                  //   input,    width = 1,                     .valid
		.snk_write_master_ready (rx_dma_write_master_response_source_ready)                   //  output,    width = 1,                     .ready
	);

	rx_dma_fifo_0 rx_dma_fifo_0 (
		.in_st_clk         (rx_dma_ftile_clock_out_clk_clk),          //   input,    width = 1,   in_st_clk.clk
		.in_st_rst         (~ftile_clk_reset_out_reset_reset),        //   input,    width = 1,   in_st_rst.reset
		.out_st_clk        (rx_dma_clock_out_clk_clk),                //   input,    width = 1,  out_st_clk.clk
		.out_st_rst        (~rx_dma_reset_out_reset_reset),           //   input,    width = 1,  out_st_rst.reset
		.csr_clk           (rx_dma_clock_out_clk_clk),                //   input,    width = 1,     csr_clk.clk
		.csr_rst           (rst_controller_001_reset_out_reset),      //   input,    width = 1,     csr_rst.reset
		.in_st_sop         (pktin_startofpacket),                     //   input,    width = 1,     in_avst.startofpacket
		.in_st_valid       (pktin_valid),                             //   input,    width = 1,            .valid
		.in_st_eop         (pktin_endofpacket),                       //   input,    width = 1,            .endofpacket
		.in_st_data        (pktin_data),                              //   input,   width = 64,            .data
		.in_st_empty       (pktin_empty),                             //   input,    width = 3,            .empty
		.in_st_error       (pktin_error),                             //   input,    width = 6,            .error
		.in_ts_valid       (rx_dma_fifo_0_in_ts_valid),               //   input,    width = 1,       in_ts.valid
		.in_ts_data        (rx_dma_fifo_0_in_ts_data),                //   input,   width = 96,            .data
		.out_st_ready      (rx_dma_fifo_0_out_avst_ready),            //   input,    width = 1,    out_avst.ready
		.out_st_sop        (rx_dma_fifo_0_out_avst_startofpacket),    //  output,    width = 1,            .startofpacket
		.out_st_valid      (rx_dma_fifo_0_out_avst_valid),            //  output,    width = 1,            .valid
		.out_st_eop        (rx_dma_fifo_0_out_avst_endofpacket),      //  output,    width = 1,            .endofpacket
		.out_st_data       (rx_dma_fifo_0_out_avst_data),             //  output,   width = 64,            .data
		.out_st_empty      (rx_dma_fifo_0_out_avst_empty),            //  output,    width = 3,            .empty
		.out_st_error      (rx_dma_fifo_0_out_avst_error),            //  output,    width = 6,            .error
		.in_ts_resp_ready  (rx_dma_dispatcher_response_source_ready), //  output,    width = 1,  in_ts_resp.ready
		.in_ts_resp_valid  (rx_dma_dispatcher_response_source_valid), //   input,    width = 1,            .valid
		.in_ts_resp_data   (rx_dma_dispatcher_response_source_data),  //   input,  width = 256,            .data
		.out_ts_resp_ready (rx_dma_fifo_0_out_ts_resp_ready),         //   input,    width = 1, out_ts_resp.ready
		.out_ts_resp_valid (rx_dma_fifo_0_out_ts_resp_valid),         //  output,    width = 1,            .valid
		.out_ts_resp_data  (rx_dma_fifo_0_out_ts_resp_data)           //  output,  width = 256,            .data
	);

	rx_dma_ftile_clock rx_dma_ftile_clock (
		.in_clk  (ftile_clk_clk),                  //   input,  width = 1,  in_clk.clk
		.out_clk (rx_dma_ftile_clock_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	rx_dma_prefetcher rx_dma_prefetcher (
		.clk                         (rx_dma_clock_out_clk_clk),                                   //   input,    width = 1,                              Clock.clk
		.reset                       (~rx_dma_reset_out_reset_reset),                              //   input,    width = 1,                        Clock_reset.reset
		.mm_read_address             (prefetcher_read_master_address),                             //  output,   width = 37,             Descriptor_Read_Master.address
		.mm_read_read                (prefetcher_read_master_read),                                //  output,    width = 1,                                   .read
		.mm_read_readdata            (prefetcher_read_master_readdata),                            //   input,  width = 128,                                   .readdata
		.mm_read_waitrequest         (prefetcher_read_master_waitrequest),                         //   input,    width = 1,                                   .waitrequest
		.mm_read_readdatavalid       (prefetcher_read_master_readdatavalid),                       //   input,    width = 1,                                   .readdatavalid
		.mm_read_burstcount          (prefetcher_read_master_burstcount),                          //  output,    width = 3,                                   .burstcount
		.mm_write_address            (prefetcher_write_master_address),                            //  output,   width = 37,            Descriptor_Write_Master.address
		.mm_write_write              (prefetcher_write_master_write),                              //  output,    width = 1,                                   .write
		.mm_write_byteenable         (prefetcher_write_master_byteenable),                         //  output,   width = 16,                                   .byteenable
		.mm_write_writedata          (prefetcher_write_master_writedata),                          //  output,  width = 128,                                   .writedata
		.mm_write_waitrequest        (prefetcher_write_master_waitrequest),                        //   input,    width = 1,                                   .waitrequest
		.mm_write_response           (prefetcher_write_master_response),                           //   input,    width = 2,                                   .response
		.mm_write_writeresponsevalid (prefetcher_write_master_writeresponsevalid),                 //   input,    width = 1,                                   .writeresponsevalid
		.st_src_descr_data           (rx_dma_prefetcher_descriptor_write_dispatcher_source_data),  //  output,  width = 256, Descriptor_Write_Dispatcher_Source.data
		.st_src_descr_valid          (rx_dma_prefetcher_descriptor_write_dispatcher_source_valid), //  output,    width = 1,                                   .valid
		.st_src_descr_ready          (rx_dma_prefetcher_descriptor_write_dispatcher_source_ready), //   input,    width = 1,                                   .ready
		.st_snk_data                 (rx_dma_fifo_0_out_ts_resp_data),                             //   input,  width = 256,                      Response_Sink.data
		.st_snk_valid                (rx_dma_fifo_0_out_ts_resp_valid),                            //   input,    width = 1,                                   .valid
		.st_snk_ready                (rx_dma_fifo_0_out_ts_resp_ready),                            //  output,    width = 1,                                   .ready
		.mm_csr_address              (mm_interconnect_0_rx_dma_prefetcher_csr_address),            //   input,    width = 3,                                Csr.address
		.mm_csr_read                 (mm_interconnect_0_rx_dma_prefetcher_csr_read),               //   input,    width = 1,                                   .read
		.mm_csr_write                (mm_interconnect_0_rx_dma_prefetcher_csr_write),              //   input,    width = 1,                                   .write
		.mm_csr_writedata            (mm_interconnect_0_rx_dma_prefetcher_csr_writedata),          //   input,   width = 32,                                   .writedata
		.mm_csr_readdata             (mm_interconnect_0_rx_dma_prefetcher_csr_readdata),           //  output,   width = 32,                                   .readdata
		.csr_irq                     (irq_irq)                                                     //  output,    width = 1,                            Csr_Irq.irq
	);

	rx_dma_reset rx_dma_reset (
		.clk         (rx_dma_clock_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_reset_n),                //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (rx_dma_reset_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	rx_dma_write_master rx_dma_write_master (
		.clk                       (rx_dma_clock_out_clk_clk),                     //   input,    width = 1,             Clock.clk
		.reset                     (~rx_dma_reset_out_reset_reset),                //   input,    width = 1,       Clock_reset.reset
		.master_address            (write_master_address),                         //  output,   width = 37, Data_Write_Master.address
		.master_write              (write_master_write),                           //  output,    width = 1,                  .write
		.master_byteenable         (write_master_byteenable),                      //  output,   width = 16,                  .byteenable
		.master_writedata          (write_master_writedata),                       //  output,  width = 128,                  .writedata
		.master_waitrequest        (write_master_waitrequest),                     //   input,    width = 1,                  .waitrequest
		.master_burstcount         (write_master_burstcount),                      //  output,    width = 5,                  .burstcount
		.master_response           (write_master_response),                        //   input,    width = 2,                  .response
		.master_writeresponsevalid (write_master_writeresponsevalid),              //   input,    width = 1,                  .writeresponsevalid
		.snk_data                  (avalon_st_adapter_out_0_data),                 //   input,  width = 128,         Data_Sink.data
		.snk_valid                 (avalon_st_adapter_out_0_valid),                //   input,    width = 1,                  .valid
		.snk_ready                 (avalon_st_adapter_out_0_ready),                //  output,    width = 1,                  .ready
		.snk_sop                   (avalon_st_adapter_out_0_startofpacket),        //   input,    width = 1,                  .startofpacket
		.snk_eop                   (avalon_st_adapter_out_0_endofpacket),          //   input,    width = 1,                  .endofpacket
		.snk_empty                 (avalon_st_adapter_out_0_empty),                //   input,    width = 4,                  .empty
		.snk_error                 (avalon_st_adapter_out_0_error),                //   input,    width = 6,                  .error
		.snk_command_data          (rx_dma_dispatcher_write_command_source_data),  //   input,  width = 256,      Command_Sink.data
		.snk_command_valid         (rx_dma_dispatcher_write_command_source_valid), //   input,    width = 1,                  .valid
		.snk_command_ready         (rx_dma_dispatcher_write_command_source_ready), //  output,    width = 1,                  .ready
		.src_response_data         (rx_dma_write_master_response_source_data),     //  output,  width = 256,   Response_Source.data
		.src_response_valid        (rx_dma_write_master_response_source_valid),    //  output,    width = 1,                  .valid
		.src_response_ready        (rx_dma_write_master_response_source_ready)     //   input,    width = 1,                  .ready
	);

	subsys_ftile_25gbe_rx_dma_altera_mm_interconnect_1920_2wjlesi mm_interconnect_0 (
		.rx_dma_csr_m0_address                                     (rx_dma_csr_m0_address),                              //   input,   width = 6,                                       rx_dma_csr_m0.address
		.rx_dma_csr_m0_waitrequest                                 (rx_dma_csr_m0_waitrequest),                          //  output,   width = 1,                                                    .waitrequest
		.rx_dma_csr_m0_burstcount                                  (rx_dma_csr_m0_burstcount),                           //   input,   width = 1,                                                    .burstcount
		.rx_dma_csr_m0_byteenable                                  (rx_dma_csr_m0_byteenable),                           //   input,   width = 4,                                                    .byteenable
		.rx_dma_csr_m0_read                                        (rx_dma_csr_m0_read),                                 //   input,   width = 1,                                                    .read
		.rx_dma_csr_m0_readdata                                    (rx_dma_csr_m0_readdata),                             //  output,  width = 32,                                                    .readdata
		.rx_dma_csr_m0_readdatavalid                               (rx_dma_csr_m0_readdatavalid),                        //  output,   width = 1,                                                    .readdatavalid
		.rx_dma_csr_m0_write                                       (rx_dma_csr_m0_write),                                //   input,   width = 1,                                                    .write
		.rx_dma_csr_m0_writedata                                   (rx_dma_csr_m0_writedata),                            //   input,  width = 32,                                                    .writedata
		.rx_dma_csr_m0_debugaccess                                 (rx_dma_csr_m0_debugaccess),                          //   input,   width = 1,                                                    .debugaccess
		.rx_dma_dispatcher_CSR_address                             (mm_interconnect_0_rx_dma_dispatcher_csr_address),    //  output,   width = 3,                               rx_dma_dispatcher_CSR.address
		.rx_dma_dispatcher_CSR_write                               (mm_interconnect_0_rx_dma_dispatcher_csr_write),      //  output,   width = 1,                                                    .write
		.rx_dma_dispatcher_CSR_read                                (mm_interconnect_0_rx_dma_dispatcher_csr_read),       //  output,   width = 1,                                                    .read
		.rx_dma_dispatcher_CSR_readdata                            (mm_interconnect_0_rx_dma_dispatcher_csr_readdata),   //   input,  width = 32,                                                    .readdata
		.rx_dma_dispatcher_CSR_writedata                           (mm_interconnect_0_rx_dma_dispatcher_csr_writedata),  //  output,  width = 32,                                                    .writedata
		.rx_dma_dispatcher_CSR_byteenable                          (mm_interconnect_0_rx_dma_dispatcher_csr_byteenable), //  output,   width = 4,                                                    .byteenable
		.rx_dma_prefetcher_Csr_address                             (mm_interconnect_0_rx_dma_prefetcher_csr_address),    //  output,   width = 3,                               rx_dma_prefetcher_Csr.address
		.rx_dma_prefetcher_Csr_write                               (mm_interconnect_0_rx_dma_prefetcher_csr_write),      //  output,   width = 1,                                                    .write
		.rx_dma_prefetcher_Csr_read                                (mm_interconnect_0_rx_dma_prefetcher_csr_read),       //  output,   width = 1,                                                    .read
		.rx_dma_prefetcher_Csr_readdata                            (mm_interconnect_0_rx_dma_prefetcher_csr_readdata),   //   input,  width = 32,                                                    .readdata
		.rx_dma_prefetcher_Csr_writedata                           (mm_interconnect_0_rx_dma_prefetcher_csr_writedata),  //  output,  width = 32,                                                    .writedata
		.rx_dma_csr_reset_reset_bridge_in_reset_reset              (~rx_dma_reset_out_reset_reset),                      //   input,   width = 1,              rx_dma_csr_reset_reset_bridge_in_reset.reset
		.rx_dma_dispatcher_clock_reset_reset_bridge_in_reset_reset (~rx_dma_reset_out_reset_reset),                      //   input,   width = 1, rx_dma_dispatcher_clock_reset_reset_bridge_in_reset.reset
		.rx_dma_clock_out_clk_clk                                  (rx_dma_clock_out_clk_clk)                            //   input,   width = 1,                                rx_dma_clock_out_clk.clk
	);

	subsys_ftile_25gbe_rx_dma_altera_avalon_st_adapter_1920_zp7psji #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (64),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (128),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (rx_dma_clock_out_clk_clk),              //   input,    width = 1, in_clk_0.clk
		.in_rst_0_reset      (~rx_dma_reset_out_reset_reset),         //   input,    width = 1, in_rst_0.reset
		.in_0_data           (rx_dma_fifo_0_out_avst_data),           //   input,   width = 64,     in_0.data
		.in_0_valid          (rx_dma_fifo_0_out_avst_valid),          //   input,    width = 1,         .valid
		.in_0_ready          (rx_dma_fifo_0_out_avst_ready),          //  output,    width = 1,         .ready
		.in_0_startofpacket  (rx_dma_fifo_0_out_avst_startofpacket),  //   input,    width = 1,         .startofpacket
		.in_0_endofpacket    (rx_dma_fifo_0_out_avst_endofpacket),    //   input,    width = 1,         .endofpacket
		.in_0_empty          (rx_dma_fifo_0_out_avst_empty),          //   input,    width = 3,         .empty
		.in_0_error          (rx_dma_fifo_0_out_avst_error),          //   input,    width = 6,         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //  output,  width = 128,    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //  output,    width = 1,         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //   input,    width = 1,         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //  output,    width = 1,         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //  output,    width = 1,         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //  output,    width = 4,         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //  output,    width = 6,         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~rx_dma_reset_out_reset_reset),  //   input,  width = 1, reset_in0.reset
		.clk            (rx_dma_ftile_clock_out_clk_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~rx_dma_reset_out_reset_reset),      //   input,  width = 1, reset_in0.reset
		.clk            (rx_dma_ftile_clock_out_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
