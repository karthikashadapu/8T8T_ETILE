// ddr4_wr_rd.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module ddr4_wr_rd (
		input  wire [20:0]  emif_mm_slave_0_address,        //     emif_mm_slave_0.address
		input  wire         emif_mm_slave_0_read,           //                    .read
		output wire [127:0] emif_mm_slave_0_readdata,       //                    .readdata
		input  wire         emif_mm_slave_0_write,          //                    .write
		input  wire [127:0] emif_mm_slave_0_writedata,      //                    .writedata
		output wire         emif_mm_slave_0_readdatavalid,  //                    .readdatavalid
		output wire         emif_mm_slave_0_waitrequest,    //                    .waitrequest
		input  wire [15:0]  emif_mm_slave_0_byteenable,     //                    .byteenable
		input  wire [6:0]   emif_mm_slave_0_burstcount,     //                    .burstcount
		input  wire         addr_span_0_cntl_read,          //    addr_span_0_cntl.read
		output wire [63:0]  addr_span_0_cntl_readdata,      //                    .readdata
		input  wire         addr_span_0_cntl_write,         //                    .write
		input  wire [63:0]  addr_span_0_cntl_writedata,     //                    .writedata
		input  wire [7:0]   addr_span_0_cntl_byteenable,    //                    .byteenable
		input  wire [20:0]  emif_mm_slave_1_address,        //     emif_mm_slave_1.address
		input  wire         emif_mm_slave_1_read,           //                    .read
		output wire [127:0] emif_mm_slave_1_readdata,       //                    .readdata
		input  wire         emif_mm_slave_1_write,          //                    .write
		input  wire [127:0] emif_mm_slave_1_writedata,      //                    .writedata
		output wire         emif_mm_slave_1_readdatavalid,  //                    .readdatavalid
		output wire         emif_mm_slave_1_waitrequest,    //                    .waitrequest
		input  wire [15:0]  emif_mm_slave_1_byteenable,     //                    .byteenable
		input  wire [6:0]   emif_mm_slave_1_burstcount,     //                    .burstcount
		input  wire         addr_span_1_cntl_read,          //    addr_span_1_cntl.read
		output wire [63:0]  addr_span_1_cntl_readdata,      //                    .readdata
		input  wire         addr_span_1_cntl_write,         //                    .write
		input  wire [63:0]  addr_span_1_cntl_writedata,     //                    .writedata
		input  wire [7:0]   addr_span_1_cntl_byteenable,    //                    .byteenable
		output wire [31:0]  wr_msgdma_ddr_address,          //       wr_msgdma_ddr.address
		output wire         wr_msgdma_ddr_read,             //                    .read
		input  wire         wr_msgdma_ddr_waitrequest,      //                    .waitrequest
		input  wire [127:0] wr_msgdma_ddr_readdata,         //                    .readdata
		output wire         wr_msgdma_ddr_write,            //                    .write
		output wire [127:0] wr_msgdma_ddr_writedata,        //                    .writedata
		input  wire         wr_msgdma_ddr_readdatavalid,    //                    .readdatavalid
		output wire [15:0]  wr_msgdma_ddr_byteenable,       //                    .byteenable
		output wire [6:0]   wr_msgdma_ddr_burstcount,       //                    .burstcount
		input  wire         in_clk_clk,                     //              in_clk.clk
		output wire         csr_bridge_s0_waitrequest,      //       csr_bridge_s0.waitrequest
		output wire [31:0]  csr_bridge_s0_readdata,         //                    .readdata
		output wire         csr_bridge_s0_readdatavalid,    //                    .readdatavalid
		input  wire [0:0]   csr_bridge_s0_burstcount,       //                    .burstcount
		input  wire [31:0]  csr_bridge_s0_writedata,        //                    .writedata
		input  wire [5:0]   csr_bridge_s0_address,          //                    .address
		input  wire         csr_bridge_s0_write,            //                    .write
		input  wire         csr_bridge_s0_read,             //                    .read
		input  wire [3:0]   csr_bridge_s0_byteenable,       //                    .byteenable
		input  wire         csr_bridge_s0_debugaccess,      //                    .debugaccess
		input  wire [12:0]  ocm_rd_address,                 //              ocm_rd.address
		input  wire         ocm_rd_read,                    //                    .read
		output wire [127:0] ocm_rd_readdata,                //                    .readdata
		input  wire         ocm_rd_clk_clk,                 //          ocm_rd_clk.clk
		input  wire         ocm_rd_reset_reset,             //        ocm_rd_reset.reset
		input  wire         ocm_rd_reset_reset_req,         //                    .reset_req
		input  wire         emif_mm_master_1_waitrequest,   //    emif_mm_master_1.waitrequest
		input  wire [127:0] emif_mm_master_1_readdata,      //                    .readdata
		input  wire         emif_mm_master_1_readdatavalid, //                    .readdatavalid
		output wire [6:0]   emif_mm_master_1_burstcount,    //                    .burstcount
		output wire [127:0] emif_mm_master_1_writedata,     //                    .writedata
		output wire [9:0]   emif_mm_master_1_address,       //                    .address
		output wire         emif_mm_master_1_write,         //                    .write
		output wire         emif_mm_master_1_read,          //                    .read
		output wire [15:0]  emif_mm_master_1_byteenable,    //                    .byteenable
		output wire         emif_mm_master_1_debugaccess,   //                    .debugaccess
		input  wire         in_reset_reset_n,               //            in_reset.reset_n
		output wire         wr_msgdma_0_csr_irq_irq,        // wr_msgdma_0_csr_irq.irq
		input  wire [127:0] wr_msgdma_0_st_sink_data,       // wr_msgdma_0_st_sink.data
		input  wire         wr_msgdma_0_st_sink_valid,      //                    .valid
		output wire         wr_msgdma_0_st_sink_ready       //                    .ready
	);

	wire          clock_bridge_0_out_clk_clk;                                             // clock_bridge_0:out_clk -> [address_span_extender_0:clk, address_span_extender_1:clk, address_span_extender_2:clk, csr_bridge:clk, intel_onchip_memory_1:clk, mm_bridge_1:clk, mm_interconnect_0:clock_bridge_0_out_clk_clk, mm_interconnect_1:clock_bridge_0_out_clk_clk, mm_interconnect_2:clock_bridge_0_out_clk_clk, reset_bridge_0:clk, rst_controller:clk, rst_controller_001:clk, wr_msgdma_0:clock_clk]
	wire          address_span_extender_1_expanded_master_waitrequest;                    // mm_interconnect_0:address_span_extender_1_expanded_master_waitrequest -> address_span_extender_1:avm_m0_waitrequest
	wire  [127:0] address_span_extender_1_expanded_master_readdata;                       // mm_interconnect_0:address_span_extender_1_expanded_master_readdata -> address_span_extender_1:avm_m0_readdata
	wire   [31:0] address_span_extender_1_expanded_master_address;                        // address_span_extender_1:avm_m0_address -> mm_interconnect_0:address_span_extender_1_expanded_master_address
	wire          address_span_extender_1_expanded_master_read;                           // address_span_extender_1:avm_m0_read -> mm_interconnect_0:address_span_extender_1_expanded_master_read
	wire   [15:0] address_span_extender_1_expanded_master_byteenable;                     // address_span_extender_1:avm_m0_byteenable -> mm_interconnect_0:address_span_extender_1_expanded_master_byteenable
	wire          address_span_extender_1_expanded_master_readdatavalid;                  // mm_interconnect_0:address_span_extender_1_expanded_master_readdatavalid -> address_span_extender_1:avm_m0_readdatavalid
	wire          address_span_extender_1_expanded_master_write;                          // address_span_extender_1:avm_m0_write -> mm_interconnect_0:address_span_extender_1_expanded_master_write
	wire  [127:0] address_span_extender_1_expanded_master_writedata;                      // address_span_extender_1:avm_m0_writedata -> mm_interconnect_0:address_span_extender_1_expanded_master_writedata
	wire    [6:0] address_span_extender_1_expanded_master_burstcount;                     // address_span_extender_1:avm_m0_burstcount -> mm_interconnect_0:address_span_extender_1_expanded_master_burstcount
	wire  [127:0] mm_interconnect_0_mm_bridge_1_s0_readdata;                              // mm_bridge_1:s0_readdata -> mm_interconnect_0:mm_bridge_1_s0_readdata
	wire          mm_interconnect_0_mm_bridge_1_s0_waitrequest;                           // mm_bridge_1:s0_waitrequest -> mm_interconnect_0:mm_bridge_1_s0_waitrequest
	wire          mm_interconnect_0_mm_bridge_1_s0_debugaccess;                           // mm_interconnect_0:mm_bridge_1_s0_debugaccess -> mm_bridge_1:s0_debugaccess
	wire    [9:0] mm_interconnect_0_mm_bridge_1_s0_address;                               // mm_interconnect_0:mm_bridge_1_s0_address -> mm_bridge_1:s0_address
	wire          mm_interconnect_0_mm_bridge_1_s0_read;                                  // mm_interconnect_0:mm_bridge_1_s0_read -> mm_bridge_1:s0_read
	wire   [15:0] mm_interconnect_0_mm_bridge_1_s0_byteenable;                            // mm_interconnect_0:mm_bridge_1_s0_byteenable -> mm_bridge_1:s0_byteenable
	wire          mm_interconnect_0_mm_bridge_1_s0_readdatavalid;                         // mm_bridge_1:s0_readdatavalid -> mm_interconnect_0:mm_bridge_1_s0_readdatavalid
	wire          mm_interconnect_0_mm_bridge_1_s0_write;                                 // mm_interconnect_0:mm_bridge_1_s0_write -> mm_bridge_1:s0_write
	wire  [127:0] mm_interconnect_0_mm_bridge_1_s0_writedata;                             // mm_interconnect_0:mm_bridge_1_s0_writedata -> mm_bridge_1:s0_writedata
	wire    [6:0] mm_interconnect_0_mm_bridge_1_s0_burstcount;                            // mm_interconnect_0:mm_bridge_1_s0_burstcount -> mm_bridge_1:s0_burstcount
	wire          csr_bridge_m0_waitrequest;                                              // mm_interconnect_1:csr_bridge_m0_waitrequest -> csr_bridge:m0_waitrequest
	wire   [31:0] csr_bridge_m0_readdata;                                                 // mm_interconnect_1:csr_bridge_m0_readdata -> csr_bridge:m0_readdata
	wire          csr_bridge_m0_debugaccess;                                              // csr_bridge:m0_debugaccess -> mm_interconnect_1:csr_bridge_m0_debugaccess
	wire    [5:0] csr_bridge_m0_address;                                                  // csr_bridge:m0_address -> mm_interconnect_1:csr_bridge_m0_address
	wire          csr_bridge_m0_read;                                                     // csr_bridge:m0_read -> mm_interconnect_1:csr_bridge_m0_read
	wire    [3:0] csr_bridge_m0_byteenable;                                               // csr_bridge:m0_byteenable -> mm_interconnect_1:csr_bridge_m0_byteenable
	wire          csr_bridge_m0_readdatavalid;                                            // mm_interconnect_1:csr_bridge_m0_readdatavalid -> csr_bridge:m0_readdatavalid
	wire   [31:0] csr_bridge_m0_writedata;                                                // csr_bridge:m0_writedata -> mm_interconnect_1:csr_bridge_m0_writedata
	wire          csr_bridge_m0_write;                                                    // csr_bridge:m0_write -> mm_interconnect_1:csr_bridge_m0_write
	wire    [0:0] csr_bridge_m0_burstcount;                                               // csr_bridge:m0_burstcount -> mm_interconnect_1:csr_bridge_m0_burstcount
	wire   [31:0] mm_interconnect_1_wr_msgdma_0_csr_readdata;                             // wr_msgdma_0:csr_readdata -> mm_interconnect_1:wr_msgdma_0_csr_readdata
	wire    [2:0] mm_interconnect_1_wr_msgdma_0_csr_address;                              // mm_interconnect_1:wr_msgdma_0_csr_address -> wr_msgdma_0:csr_address
	wire          mm_interconnect_1_wr_msgdma_0_csr_read;                                 // mm_interconnect_1:wr_msgdma_0_csr_read -> wr_msgdma_0:csr_read
	wire    [3:0] mm_interconnect_1_wr_msgdma_0_csr_byteenable;                           // mm_interconnect_1:wr_msgdma_0_csr_byteenable -> wr_msgdma_0:csr_byteenable
	wire          mm_interconnect_1_wr_msgdma_0_csr_write;                                // mm_interconnect_1:wr_msgdma_0_csr_write -> wr_msgdma_0:csr_write
	wire   [31:0] mm_interconnect_1_wr_msgdma_0_csr_writedata;                            // mm_interconnect_1:wr_msgdma_0_csr_writedata -> wr_msgdma_0:csr_writedata
	wire          mm_interconnect_1_wr_msgdma_0_descriptor_slave_waitrequest;             // wr_msgdma_0:descriptor_slave_waitrequest -> mm_interconnect_1:wr_msgdma_0_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_1_wr_msgdma_0_descriptor_slave_byteenable;              // mm_interconnect_1:wr_msgdma_0_descriptor_slave_byteenable -> wr_msgdma_0:descriptor_slave_byteenable
	wire          mm_interconnect_1_wr_msgdma_0_descriptor_slave_write;                   // mm_interconnect_1:wr_msgdma_0_descriptor_slave_write -> wr_msgdma_0:descriptor_slave_write
	wire  [127:0] mm_interconnect_1_wr_msgdma_0_descriptor_slave_writedata;               // mm_interconnect_1:wr_msgdma_0_descriptor_slave_writedata -> wr_msgdma_0:descriptor_slave_writedata
	wire          wr_msgdma_0_mm_write_waitrequest;                                       // mm_interconnect_2:wr_msgdma_0_mm_write_waitrequest -> wr_msgdma_0:mm_write_waitrequest
	wire   [31:0] wr_msgdma_0_mm_write_address;                                           // wr_msgdma_0:mm_write_address -> mm_interconnect_2:wr_msgdma_0_mm_write_address
	wire   [15:0] wr_msgdma_0_mm_write_byteenable;                                        // wr_msgdma_0:mm_write_byteenable -> mm_interconnect_2:wr_msgdma_0_mm_write_byteenable
	wire          wr_msgdma_0_mm_write_write;                                             // wr_msgdma_0:mm_write_write -> mm_interconnect_2:wr_msgdma_0_mm_write_write
	wire  [127:0] wr_msgdma_0_mm_write_writedata;                                         // wr_msgdma_0:mm_write_writedata -> mm_interconnect_2:wr_msgdma_0_mm_write_writedata
	wire    [6:0] wr_msgdma_0_mm_write_burstcount;                                        // wr_msgdma_0:mm_write_burstcount -> mm_interconnect_2:wr_msgdma_0_mm_write_burstcount
	wire   [12:0] mm_interconnect_2_intel_onchip_memory_1_s1_address;                     // mm_interconnect_2:intel_onchip_memory_1_s1_address -> intel_onchip_memory_1:address
	wire   [15:0] mm_interconnect_2_intel_onchip_memory_1_s1_byteenable;                  // mm_interconnect_2:intel_onchip_memory_1_s1_byteenable -> intel_onchip_memory_1:byteenable
	wire          mm_interconnect_2_intel_onchip_memory_1_s1_write;                       // mm_interconnect_2:intel_onchip_memory_1_s1_write -> intel_onchip_memory_1:write
	wire  [127:0] mm_interconnect_2_intel_onchip_memory_1_s1_writedata;                   // mm_interconnect_2:intel_onchip_memory_1_s1_writedata -> intel_onchip_memory_1:writedata
	wire  [127:0] mm_interconnect_2_address_span_extender_2_windowed_slave_readdata;      // address_span_extender_2:avs_s0_readdata -> mm_interconnect_2:address_span_extender_2_windowed_slave_readdata
	wire          mm_interconnect_2_address_span_extender_2_windowed_slave_waitrequest;   // address_span_extender_2:avs_s0_waitrequest -> mm_interconnect_2:address_span_extender_2_windowed_slave_waitrequest
	wire   [20:0] mm_interconnect_2_address_span_extender_2_windowed_slave_address;       // mm_interconnect_2:address_span_extender_2_windowed_slave_address -> address_span_extender_2:avs_s0_address
	wire          mm_interconnect_2_address_span_extender_2_windowed_slave_read;          // mm_interconnect_2:address_span_extender_2_windowed_slave_read -> address_span_extender_2:avs_s0_read
	wire   [15:0] mm_interconnect_2_address_span_extender_2_windowed_slave_byteenable;    // mm_interconnect_2:address_span_extender_2_windowed_slave_byteenable -> address_span_extender_2:avs_s0_byteenable
	wire          mm_interconnect_2_address_span_extender_2_windowed_slave_readdatavalid; // address_span_extender_2:avs_s0_readdatavalid -> mm_interconnect_2:address_span_extender_2_windowed_slave_readdatavalid
	wire          mm_interconnect_2_address_span_extender_2_windowed_slave_write;         // mm_interconnect_2:address_span_extender_2_windowed_slave_write -> address_span_extender_2:avs_s0_write
	wire  [127:0] mm_interconnect_2_address_span_extender_2_windowed_slave_writedata;     // mm_interconnect_2:address_span_extender_2_windowed_slave_writedata -> address_span_extender_2:avs_s0_writedata
	wire    [6:0] mm_interconnect_2_address_span_extender_2_windowed_slave_burstcount;    // mm_interconnect_2:address_span_extender_2_windowed_slave_burstcount -> address_span_extender_2:avs_s0_burstcount
	wire          rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [address_span_extender_0:reset, address_span_extender_1:reset, address_span_extender_2:reset, csr_bridge:reset, intel_onchip_memory_1:reset, mm_bridge_1:reset, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                                     // rst_controller:reset_req -> [intel_onchip_memory_1:reset_req, rst_translator:reset_req_in]
	wire          reset_bridge_0_out_reset_reset;                                         // reset_bridge_0:out_reset_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                     // rst_controller_001:reset_out -> [mm_interconnect_0:address_span_extender_1_expanded_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:csr_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:wr_msgdma_0_reset_n_reset_bridge_in_reset_reset, mm_interconnect_2:intel_onchip_memory_1_reset1_reset_bridge_in_reset_reset, mm_interconnect_2:wr_msgdma_0_reset_n_reset_bridge_in_reset_reset, wr_msgdma_0:reset_n_reset_n]

	ed_synth_address_span_extender_0 address_span_extender_0 (
		.clk                  (clock_bridge_0_out_clk_clk),     //   input,    width = 1,           clock.clk
		.reset                (rst_controller_reset_out_reset), //   input,    width = 1,           reset.reset
		.avs_s0_address       (emif_mm_slave_0_address),        //   input,   width = 21,  windowed_slave.address
		.avs_s0_read          (emif_mm_slave_0_read),           //   input,    width = 1,                .read
		.avs_s0_readdata      (emif_mm_slave_0_readdata),       //  output,  width = 128,                .readdata
		.avs_s0_write         (emif_mm_slave_0_write),          //   input,    width = 1,                .write
		.avs_s0_writedata     (emif_mm_slave_0_writedata),      //   input,  width = 128,                .writedata
		.avs_s0_readdatavalid (emif_mm_slave_0_readdatavalid),  //  output,    width = 1,                .readdatavalid
		.avs_s0_waitrequest   (emif_mm_slave_0_waitrequest),    //  output,    width = 1,                .waitrequest
		.avs_s0_byteenable    (emif_mm_slave_0_byteenable),     //   input,   width = 16,                .byteenable
		.avs_s0_burstcount    (emif_mm_slave_0_burstcount),     //   input,    width = 7,                .burstcount
		.avm_m0_address       (),                               //  output,   width = 32, expanded_master.address
		.avm_m0_read          (),                               //  output,    width = 1,                .read
		.avm_m0_waitrequest   (),                               //   input,    width = 1,                .waitrequest
		.avm_m0_readdata      (),                               //   input,  width = 128,                .readdata
		.avm_m0_write         (),                               //  output,    width = 1,                .write
		.avm_m0_writedata     (),                               //  output,  width = 128,                .writedata
		.avm_m0_readdatavalid (),                               //   input,    width = 1,                .readdatavalid
		.avm_m0_byteenable    (),                               //  output,   width = 16,                .byteenable
		.avm_m0_burstcount    (),                               //  output,    width = 7,                .burstcount
		.avs_cntl_read        (addr_span_0_cntl_read),          //   input,    width = 1,            cntl.read
		.avs_cntl_readdata    (addr_span_0_cntl_readdata),      //  output,   width = 64,                .readdata
		.avs_cntl_write       (addr_span_0_cntl_write),         //   input,    width = 1,                .write
		.avs_cntl_writedata   (addr_span_0_cntl_writedata),     //   input,   width = 64,                .writedata
		.avs_cntl_byteenable  (addr_span_0_cntl_byteenable)     //   input,    width = 8,                .byteenable
	);

	ed_synth_address_span_extender_0 address_span_extender_1 (
		.clk                  (clock_bridge_0_out_clk_clk),                            //   input,    width = 1,           clock.clk
		.reset                (rst_controller_reset_out_reset),                        //   input,    width = 1,           reset.reset
		.avs_s0_address       (emif_mm_slave_1_address),                               //   input,   width = 21,  windowed_slave.address
		.avs_s0_read          (emif_mm_slave_1_read),                                  //   input,    width = 1,                .read
		.avs_s0_readdata      (emif_mm_slave_1_readdata),                              //  output,  width = 128,                .readdata
		.avs_s0_write         (emif_mm_slave_1_write),                                 //   input,    width = 1,                .write
		.avs_s0_writedata     (emif_mm_slave_1_writedata),                             //   input,  width = 128,                .writedata
		.avs_s0_readdatavalid (emif_mm_slave_1_readdatavalid),                         //  output,    width = 1,                .readdatavalid
		.avs_s0_waitrequest   (emif_mm_slave_1_waitrequest),                           //  output,    width = 1,                .waitrequest
		.avs_s0_byteenable    (emif_mm_slave_1_byteenable),                            //   input,   width = 16,                .byteenable
		.avs_s0_burstcount    (emif_mm_slave_1_burstcount),                            //   input,    width = 7,                .burstcount
		.avm_m0_address       (address_span_extender_1_expanded_master_address),       //  output,   width = 32, expanded_master.address
		.avm_m0_read          (address_span_extender_1_expanded_master_read),          //  output,    width = 1,                .read
		.avm_m0_waitrequest   (address_span_extender_1_expanded_master_waitrequest),   //   input,    width = 1,                .waitrequest
		.avm_m0_readdata      (address_span_extender_1_expanded_master_readdata),      //   input,  width = 128,                .readdata
		.avm_m0_write         (address_span_extender_1_expanded_master_write),         //  output,    width = 1,                .write
		.avm_m0_writedata     (address_span_extender_1_expanded_master_writedata),     //  output,  width = 128,                .writedata
		.avm_m0_readdatavalid (address_span_extender_1_expanded_master_readdatavalid), //   input,    width = 1,                .readdatavalid
		.avm_m0_byteenable    (address_span_extender_1_expanded_master_byteenable),    //  output,   width = 16,                .byteenable
		.avm_m0_burstcount    (address_span_extender_1_expanded_master_burstcount),    //  output,    width = 7,                .burstcount
		.avs_cntl_read        (addr_span_1_cntl_read),                                 //   input,    width = 1,            cntl.read
		.avs_cntl_readdata    (addr_span_1_cntl_readdata),                             //  output,   width = 64,                .readdata
		.avs_cntl_write       (addr_span_1_cntl_write),                                //   input,    width = 1,                .write
		.avs_cntl_writedata   (addr_span_1_cntl_writedata),                            //   input,   width = 64,                .writedata
		.avs_cntl_byteenable  (addr_span_1_cntl_byteenable)                            //   input,    width = 8,                .byteenable
	);

	ddr4_wr_rd_address_span_extender_2 address_span_extender_2 (
		.clk                  (clock_bridge_0_out_clk_clk),                                             //   input,    width = 1,           clock.clk
		.reset                (rst_controller_reset_out_reset),                                         //   input,    width = 1,           reset.reset
		.avs_s0_address       (mm_interconnect_2_address_span_extender_2_windowed_slave_address),       //   input,   width = 21,  windowed_slave.address
		.avs_s0_read          (mm_interconnect_2_address_span_extender_2_windowed_slave_read),          //   input,    width = 1,                .read
		.avs_s0_readdata      (mm_interconnect_2_address_span_extender_2_windowed_slave_readdata),      //  output,  width = 128,                .readdata
		.avs_s0_write         (mm_interconnect_2_address_span_extender_2_windowed_slave_write),         //   input,    width = 1,                .write
		.avs_s0_writedata     (mm_interconnect_2_address_span_extender_2_windowed_slave_writedata),     //   input,  width = 128,                .writedata
		.avs_s0_readdatavalid (mm_interconnect_2_address_span_extender_2_windowed_slave_readdatavalid), //  output,    width = 1,                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_2_address_span_extender_2_windowed_slave_waitrequest),   //  output,    width = 1,                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_2_address_span_extender_2_windowed_slave_byteenable),    //   input,   width = 16,                .byteenable
		.avs_s0_burstcount    (mm_interconnect_2_address_span_extender_2_windowed_slave_burstcount),    //   input,    width = 7,                .burstcount
		.avm_m0_address       (wr_msgdma_ddr_address),                                                  //  output,   width = 32, expanded_master.address
		.avm_m0_read          (wr_msgdma_ddr_read),                                                     //  output,    width = 1,                .read
		.avm_m0_waitrequest   (wr_msgdma_ddr_waitrequest),                                              //   input,    width = 1,                .waitrequest
		.avm_m0_readdata      (wr_msgdma_ddr_readdata),                                                 //   input,  width = 128,                .readdata
		.avm_m0_write         (wr_msgdma_ddr_write),                                                    //  output,    width = 1,                .write
		.avm_m0_writedata     (wr_msgdma_ddr_writedata),                                                //  output,  width = 128,                .writedata
		.avm_m0_readdatavalid (wr_msgdma_ddr_readdatavalid),                                            //   input,    width = 1,                .readdatavalid
		.avm_m0_byteenable    (wr_msgdma_ddr_byteenable),                                               //  output,   width = 16,                .byteenable
		.avm_m0_burstcount    (wr_msgdma_ddr_burstcount),                                               //  output,    width = 7,                .burstcount
		.avs_cntl_read        (),                                                                       //   input,    width = 1,            cntl.read
		.avs_cntl_readdata    (),                                                                       //  output,   width = 64,                .readdata
		.avs_cntl_write       (),                                                                       //   input,    width = 1,                .write
		.avs_cntl_writedata   (),                                                                       //   input,   width = 64,                .writedata
		.avs_cntl_byteenable  ()                                                                        //   input,    width = 8,                .byteenable
	);

	ddr4_wr_rd_clock_bridge_0 clock_bridge_0 (
		.in_clk  (in_clk_clk),                 //   input,  width = 1,  in_clk.clk
		.out_clk (clock_bridge_0_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	ddr4_wr_rd_mm_bridge_1 csr_bridge (
		.clk              (clock_bridge_0_out_clk_clk),     //   input,   width = 1,   clk.clk
		.reset            (rst_controller_reset_out_reset), //   input,   width = 1, reset.reset
		.s0_waitrequest   (csr_bridge_s0_waitrequest),      //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (csr_bridge_s0_readdata),         //  output,  width = 32,      .readdata
		.s0_readdatavalid (csr_bridge_s0_readdatavalid),    //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (csr_bridge_s0_burstcount),       //   input,   width = 1,      .burstcount
		.s0_writedata     (csr_bridge_s0_writedata),        //   input,  width = 32,      .writedata
		.s0_address       (csr_bridge_s0_address),          //   input,   width = 6,      .address
		.s0_write         (csr_bridge_s0_write),            //   input,   width = 1,      .write
		.s0_read          (csr_bridge_s0_read),             //   input,   width = 1,      .read
		.s0_byteenable    (csr_bridge_s0_byteenable),       //   input,   width = 4,      .byteenable
		.s0_debugaccess   (csr_bridge_s0_debugaccess),      //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (csr_bridge_m0_waitrequest),      //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (csr_bridge_m0_readdata),         //   input,  width = 32,      .readdata
		.m0_readdatavalid (csr_bridge_m0_readdatavalid),    //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (csr_bridge_m0_burstcount),       //  output,   width = 1,      .burstcount
		.m0_writedata     (csr_bridge_m0_writedata),        //  output,  width = 32,      .writedata
		.m0_address       (csr_bridge_m0_address),          //  output,   width = 6,      .address
		.m0_write         (csr_bridge_m0_write),            //  output,   width = 1,      .write
		.m0_read          (csr_bridge_m0_read),             //  output,   width = 1,      .read
		.m0_byteenable    (csr_bridge_m0_byteenable),       //  output,   width = 4,      .byteenable
		.m0_debugaccess   (csr_bridge_m0_debugaccess)       //  output,   width = 1,      .debugaccess
	);

	ddr4_wr_rd_intel_onchip_memory_1 intel_onchip_memory_1 (
		.clk        (clock_bridge_0_out_clk_clk),                            //   input,    width = 1,   clk1.clk
		.address    (mm_interconnect_2_intel_onchip_memory_1_s1_address),    //   input,   width = 13,     s1.address
		.byteenable (mm_interconnect_2_intel_onchip_memory_1_s1_byteenable), //   input,   width = 16,       .byteenable
		.write      (mm_interconnect_2_intel_onchip_memory_1_s1_write),      //   input,    width = 1,       .write
		.writedata  (mm_interconnect_2_intel_onchip_memory_1_s1_writedata),  //   input,  width = 128,       .writedata
		.reset      (rst_controller_reset_out_reset),                        //   input,    width = 1, reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                    //   input,    width = 1,       .reset_req
		.address2   (ocm_rd_address),                                        //   input,   width = 13,     s2.address
		.read2      (ocm_rd_read),                                           //   input,    width = 1,       .read
		.readdata2  (ocm_rd_readdata),                                       //  output,  width = 128,       .readdata
		.clk2       (ocm_rd_clk_clk),                                        //   input,    width = 1,   clk2.clk
		.reset2     (ocm_rd_reset_reset),                                    //   input,    width = 1, reset2.reset
		.reset_req2 (ocm_rd_reset_reset_req)                                 //   input,    width = 1,       .reset_req
	);

	ed_synth_mm_bridge_0 mm_bridge_1 (
		.clk              (clock_bridge_0_out_clk_clk),                     //   input,    width = 1,   clk.clk
		.reset            (rst_controller_reset_out_reset),                 //   input,    width = 1, reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_1_s0_waitrequest),   //  output,    width = 1,    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_1_s0_readdata),      //  output,  width = 128,      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_1_s0_readdatavalid), //  output,    width = 1,      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_1_s0_burstcount),    //   input,    width = 7,      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_1_s0_writedata),     //   input,  width = 128,      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_1_s0_address),       //   input,   width = 10,      .address
		.s0_write         (mm_interconnect_0_mm_bridge_1_s0_write),         //   input,    width = 1,      .write
		.s0_read          (mm_interconnect_0_mm_bridge_1_s0_read),          //   input,    width = 1,      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_1_s0_byteenable),    //   input,   width = 16,      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_1_s0_debugaccess),   //   input,    width = 1,      .debugaccess
		.m0_waitrequest   (emif_mm_master_1_waitrequest),                   //   input,    width = 1,    m0.waitrequest
		.m0_readdata      (emif_mm_master_1_readdata),                      //   input,  width = 128,      .readdata
		.m0_readdatavalid (emif_mm_master_1_readdatavalid),                 //   input,    width = 1,      .readdatavalid
		.m0_burstcount    (emif_mm_master_1_burstcount),                    //  output,    width = 7,      .burstcount
		.m0_writedata     (emif_mm_master_1_writedata),                     //  output,  width = 128,      .writedata
		.m0_address       (emif_mm_master_1_address),                       //  output,   width = 10,      .address
		.m0_write         (emif_mm_master_1_write),                         //  output,    width = 1,      .write
		.m0_read          (emif_mm_master_1_read),                          //  output,    width = 1,      .read
		.m0_byteenable    (emif_mm_master_1_byteenable),                    //  output,   width = 16,      .byteenable
		.m0_debugaccess   (emif_mm_master_1_debugaccess)                    //  output,    width = 1,      .debugaccess
	);

	ddr4_wr_rd_reset_bridge_0 reset_bridge_0 (
		.clk         (clock_bridge_0_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (in_reset_reset_n),               //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (reset_bridge_0_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	ed_synth_msgdma_0 wr_msgdma_0 (
		.clock_clk                    (clock_bridge_0_out_clk_clk),                                 //   input,    width = 1,            clock.clk
		.reset_n_reset_n              (~rst_controller_001_reset_out_reset),                        //   input,    width = 1,          reset_n.reset_n
		.csr_writedata                (mm_interconnect_1_wr_msgdma_0_csr_writedata),                //   input,   width = 32,              csr.writedata
		.csr_write                    (mm_interconnect_1_wr_msgdma_0_csr_write),                    //   input,    width = 1,                 .write
		.csr_byteenable               (mm_interconnect_1_wr_msgdma_0_csr_byteenable),               //   input,    width = 4,                 .byteenable
		.csr_readdata                 (mm_interconnect_1_wr_msgdma_0_csr_readdata),                 //  output,   width = 32,                 .readdata
		.csr_read                     (mm_interconnect_1_wr_msgdma_0_csr_read),                     //   input,    width = 1,                 .read
		.csr_address                  (mm_interconnect_1_wr_msgdma_0_csr_address),                  //   input,    width = 3,                 .address
		.descriptor_slave_write       (mm_interconnect_1_wr_msgdma_0_descriptor_slave_write),       //   input,    width = 1, descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_1_wr_msgdma_0_descriptor_slave_waitrequest), //  output,    width = 1,                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_1_wr_msgdma_0_descriptor_slave_writedata),   //   input,  width = 128,                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_1_wr_msgdma_0_descriptor_slave_byteenable),  //   input,   width = 16,                 .byteenable
		.csr_irq_irq                  (wr_msgdma_0_csr_irq_irq),                                    //  output,    width = 1,          csr_irq.irq
		.mm_write_address             (wr_msgdma_0_mm_write_address),                               //  output,   width = 32,         mm_write.address
		.mm_write_write               (wr_msgdma_0_mm_write_write),                                 //  output,    width = 1,                 .write
		.mm_write_byteenable          (wr_msgdma_0_mm_write_byteenable),                            //  output,   width = 16,                 .byteenable
		.mm_write_writedata           (wr_msgdma_0_mm_write_writedata),                             //  output,  width = 128,                 .writedata
		.mm_write_waitrequest         (wr_msgdma_0_mm_write_waitrequest),                           //   input,    width = 1,                 .waitrequest
		.mm_write_burstcount          (wr_msgdma_0_mm_write_burstcount),                            //  output,    width = 7,                 .burstcount
		.st_sink_data                 (wr_msgdma_0_st_sink_data),                                   //   input,  width = 128,          st_sink.data
		.st_sink_valid                (wr_msgdma_0_st_sink_valid),                                  //   input,    width = 1,                 .valid
		.st_sink_ready                (wr_msgdma_0_st_sink_ready)                                   //  output,    width = 1,                 .ready
	);

	ddr4_wr_rd_altera_mm_interconnect_1920_co3wyjy mm_interconnect_0 (
		.address_span_extender_1_expanded_master_address                                      (address_span_extender_1_expanded_master_address),       //   input,   width = 32,                                        address_span_extender_1_expanded_master.address
		.address_span_extender_1_expanded_master_waitrequest                                  (address_span_extender_1_expanded_master_waitrequest),   //  output,    width = 1,                                                                               .waitrequest
		.address_span_extender_1_expanded_master_burstcount                                   (address_span_extender_1_expanded_master_burstcount),    //   input,    width = 7,                                                                               .burstcount
		.address_span_extender_1_expanded_master_byteenable                                   (address_span_extender_1_expanded_master_byteenable),    //   input,   width = 16,                                                                               .byteenable
		.address_span_extender_1_expanded_master_read                                         (address_span_extender_1_expanded_master_read),          //   input,    width = 1,                                                                               .read
		.address_span_extender_1_expanded_master_readdata                                     (address_span_extender_1_expanded_master_readdata),      //  output,  width = 128,                                                                               .readdata
		.address_span_extender_1_expanded_master_readdatavalid                                (address_span_extender_1_expanded_master_readdatavalid), //  output,    width = 1,                                                                               .readdatavalid
		.address_span_extender_1_expanded_master_write                                        (address_span_extender_1_expanded_master_write),         //   input,    width = 1,                                                                               .write
		.address_span_extender_1_expanded_master_writedata                                    (address_span_extender_1_expanded_master_writedata),     //   input,  width = 128,                                                                               .writedata
		.mm_bridge_1_s0_address                                                               (mm_interconnect_0_mm_bridge_1_s0_address),              //  output,   width = 10,                                                                 mm_bridge_1_s0.address
		.mm_bridge_1_s0_write                                                                 (mm_interconnect_0_mm_bridge_1_s0_write),                //  output,    width = 1,                                                                               .write
		.mm_bridge_1_s0_read                                                                  (mm_interconnect_0_mm_bridge_1_s0_read),                 //  output,    width = 1,                                                                               .read
		.mm_bridge_1_s0_readdata                                                              (mm_interconnect_0_mm_bridge_1_s0_readdata),             //   input,  width = 128,                                                                               .readdata
		.mm_bridge_1_s0_writedata                                                             (mm_interconnect_0_mm_bridge_1_s0_writedata),            //  output,  width = 128,                                                                               .writedata
		.mm_bridge_1_s0_burstcount                                                            (mm_interconnect_0_mm_bridge_1_s0_burstcount),           //  output,    width = 7,                                                                               .burstcount
		.mm_bridge_1_s0_byteenable                                                            (mm_interconnect_0_mm_bridge_1_s0_byteenable),           //  output,   width = 16,                                                                               .byteenable
		.mm_bridge_1_s0_readdatavalid                                                         (mm_interconnect_0_mm_bridge_1_s0_readdatavalid),        //   input,    width = 1,                                                                               .readdatavalid
		.mm_bridge_1_s0_waitrequest                                                           (mm_interconnect_0_mm_bridge_1_s0_waitrequest),          //   input,    width = 1,                                                                               .waitrequest
		.mm_bridge_1_s0_debugaccess                                                           (mm_interconnect_0_mm_bridge_1_s0_debugaccess),          //  output,    width = 1,                                                                               .debugaccess
		.address_span_extender_1_expanded_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    //   input,    width = 1, address_span_extender_1_expanded_master_translator_reset_reset_bridge_in_reset.reset
		.clock_bridge_0_out_clk_clk                                                           (clock_bridge_0_out_clk_clk)                             //   input,    width = 1,                                                         clock_bridge_0_out_clk.clk
	);

	ddr4_wr_rd_altera_mm_interconnect_1920_dgurhwa mm_interconnect_1 (
		.csr_bridge_m0_address                           (csr_bridge_m0_address),                                      //   input,    width = 6,                             csr_bridge_m0.address
		.csr_bridge_m0_waitrequest                       (csr_bridge_m0_waitrequest),                                  //  output,    width = 1,                                          .waitrequest
		.csr_bridge_m0_burstcount                        (csr_bridge_m0_burstcount),                                   //   input,    width = 1,                                          .burstcount
		.csr_bridge_m0_byteenable                        (csr_bridge_m0_byteenable),                                   //   input,    width = 4,                                          .byteenable
		.csr_bridge_m0_read                              (csr_bridge_m0_read),                                         //   input,    width = 1,                                          .read
		.csr_bridge_m0_readdata                          (csr_bridge_m0_readdata),                                     //  output,   width = 32,                                          .readdata
		.csr_bridge_m0_readdatavalid                     (csr_bridge_m0_readdatavalid),                                //  output,    width = 1,                                          .readdatavalid
		.csr_bridge_m0_write                             (csr_bridge_m0_write),                                        //   input,    width = 1,                                          .write
		.csr_bridge_m0_writedata                         (csr_bridge_m0_writedata),                                    //   input,   width = 32,                                          .writedata
		.csr_bridge_m0_debugaccess                       (csr_bridge_m0_debugaccess),                                  //   input,    width = 1,                                          .debugaccess
		.wr_msgdma_0_csr_address                         (mm_interconnect_1_wr_msgdma_0_csr_address),                  //  output,    width = 3,                           wr_msgdma_0_csr.address
		.wr_msgdma_0_csr_write                           (mm_interconnect_1_wr_msgdma_0_csr_write),                    //  output,    width = 1,                                          .write
		.wr_msgdma_0_csr_read                            (mm_interconnect_1_wr_msgdma_0_csr_read),                     //  output,    width = 1,                                          .read
		.wr_msgdma_0_csr_readdata                        (mm_interconnect_1_wr_msgdma_0_csr_readdata),                 //   input,   width = 32,                                          .readdata
		.wr_msgdma_0_csr_writedata                       (mm_interconnect_1_wr_msgdma_0_csr_writedata),                //  output,   width = 32,                                          .writedata
		.wr_msgdma_0_csr_byteenable                      (mm_interconnect_1_wr_msgdma_0_csr_byteenable),               //  output,    width = 4,                                          .byteenable
		.wr_msgdma_0_descriptor_slave_write              (mm_interconnect_1_wr_msgdma_0_descriptor_slave_write),       //  output,    width = 1,              wr_msgdma_0_descriptor_slave.write
		.wr_msgdma_0_descriptor_slave_writedata          (mm_interconnect_1_wr_msgdma_0_descriptor_slave_writedata),   //  output,  width = 128,                                          .writedata
		.wr_msgdma_0_descriptor_slave_byteenable         (mm_interconnect_1_wr_msgdma_0_descriptor_slave_byteenable),  //  output,   width = 16,                                          .byteenable
		.wr_msgdma_0_descriptor_slave_waitrequest        (mm_interconnect_1_wr_msgdma_0_descriptor_slave_waitrequest), //   input,    width = 1,                                          .waitrequest
		.csr_bridge_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                         //   input,    width = 1,    csr_bridge_reset_reset_bridge_in_reset.reset
		.wr_msgdma_0_reset_n_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         //   input,    width = 1, wr_msgdma_0_reset_n_reset_bridge_in_reset.reset
		.clock_bridge_0_out_clk_clk                      (clock_bridge_0_out_clk_clk)                                  //   input,    width = 1,                    clock_bridge_0_out_clk.clk
	);

	ddr4_wr_rd_altera_mm_interconnect_1920_6lb3vry mm_interconnect_2 (
		.wr_msgdma_0_mm_write_address                             (wr_msgdma_0_mm_write_address),                                           //   input,   width = 32,                               wr_msgdma_0_mm_write.address
		.wr_msgdma_0_mm_write_waitrequest                         (wr_msgdma_0_mm_write_waitrequest),                                       //  output,    width = 1,                                                   .waitrequest
		.wr_msgdma_0_mm_write_burstcount                          (wr_msgdma_0_mm_write_burstcount),                                        //   input,    width = 7,                                                   .burstcount
		.wr_msgdma_0_mm_write_byteenable                          (wr_msgdma_0_mm_write_byteenable),                                        //   input,   width = 16,                                                   .byteenable
		.wr_msgdma_0_mm_write_write                               (wr_msgdma_0_mm_write_write),                                             //   input,    width = 1,                                                   .write
		.wr_msgdma_0_mm_write_writedata                           (wr_msgdma_0_mm_write_writedata),                                         //   input,  width = 128,                                                   .writedata
		.intel_onchip_memory_1_s1_address                         (mm_interconnect_2_intel_onchip_memory_1_s1_address),                     //  output,   width = 13,                           intel_onchip_memory_1_s1.address
		.intel_onchip_memory_1_s1_write                           (mm_interconnect_2_intel_onchip_memory_1_s1_write),                       //  output,    width = 1,                                                   .write
		.intel_onchip_memory_1_s1_writedata                       (mm_interconnect_2_intel_onchip_memory_1_s1_writedata),                   //  output,  width = 128,                                                   .writedata
		.intel_onchip_memory_1_s1_byteenable                      (mm_interconnect_2_intel_onchip_memory_1_s1_byteenable),                  //  output,   width = 16,                                                   .byteenable
		.address_span_extender_2_windowed_slave_address           (mm_interconnect_2_address_span_extender_2_windowed_slave_address),       //  output,   width = 21,             address_span_extender_2_windowed_slave.address
		.address_span_extender_2_windowed_slave_write             (mm_interconnect_2_address_span_extender_2_windowed_slave_write),         //  output,    width = 1,                                                   .write
		.address_span_extender_2_windowed_slave_read              (mm_interconnect_2_address_span_extender_2_windowed_slave_read),          //  output,    width = 1,                                                   .read
		.address_span_extender_2_windowed_slave_readdata          (mm_interconnect_2_address_span_extender_2_windowed_slave_readdata),      //   input,  width = 128,                                                   .readdata
		.address_span_extender_2_windowed_slave_writedata         (mm_interconnect_2_address_span_extender_2_windowed_slave_writedata),     //  output,  width = 128,                                                   .writedata
		.address_span_extender_2_windowed_slave_burstcount        (mm_interconnect_2_address_span_extender_2_windowed_slave_burstcount),    //  output,    width = 7,                                                   .burstcount
		.address_span_extender_2_windowed_slave_byteenable        (mm_interconnect_2_address_span_extender_2_windowed_slave_byteenable),    //  output,   width = 16,                                                   .byteenable
		.address_span_extender_2_windowed_slave_readdatavalid     (mm_interconnect_2_address_span_extender_2_windowed_slave_readdatavalid), //   input,    width = 1,                                                   .readdatavalid
		.address_span_extender_2_windowed_slave_waitrequest       (mm_interconnect_2_address_span_extender_2_windowed_slave_waitrequest),   //   input,    width = 1,                                                   .waitrequest
		.wr_msgdma_0_reset_n_reset_bridge_in_reset_reset          (rst_controller_001_reset_out_reset),                                     //   input,    width = 1,          wr_msgdma_0_reset_n_reset_bridge_in_reset.reset
		.intel_onchip_memory_1_reset1_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                     //   input,    width = 1, intel_onchip_memory_1_reset1_reset_bridge_in_reset.reset
		.clock_bridge_0_out_clk_clk                               (clock_bridge_0_out_clk_clk)                                              //   input,    width = 1,                             clock_bridge_0_out_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_bridge_0_out_reset_reset),    //   input,  width = 1, reset_in0.reset
		.clk            (clock_bridge_0_out_clk_clk),         //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_bridge_0_out_reset_reset),    //   input,  width = 1, reset_in0.reset
		.clk            (clock_bridge_0_out_clk_clk),         //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
