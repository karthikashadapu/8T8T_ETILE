// subsys_ftile_25gbe_tx_dma.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module subsys_ftile_25gbe_tx_dma #(
		parameter FP_WIDTH = 8
	) (
		input  wire [0:0]   ts_chs_compl_0_clk_bus_in_clk,              // ts_chs_compl_0_clk_bus_in.clk
		input  wire [0:0]   ts_chs_compl_0_rst_bus_in_reset,            // ts_chs_compl_0_rst_bus_in.reset
		input  wire [0:0]   ts_chs_compl_0_i_ts_valid,                  //       ts_chs_compl_0_i_ts.valid
		input  wire [19:0]  ts_chs_compl_0_i_ts_fingerprint,            //                          .fingerprint
		input  wire [95:0]  ts_chs_compl_0_i_ts_data,                   //                          .data
		input  wire         dma_clk_clk,                                //                   dma_clk.clk
		output wire         csr_waitrequest,                            //                       csr.waitrequest
		output wire [31:0]  csr_readdata,                               //                          .readdata
		output wire         csr_readdatavalid,                          //                          .readdatavalid
		input  wire [0:0]   csr_burstcount,                             //                          .burstcount
		input  wire [31:0]  csr_writedata,                              //                          .writedata
		input  wire [5:0]   csr_address,                                //                          .address
		input  wire         csr_write,                                  //                          .write
		input  wire         csr_read,                                   //                          .read
		input  wire [3:0]   csr_byteenable,                             //                          .byteenable
		input  wire         csr_debugaccess,                            //                          .debugaccess
		input  wire         tx_dma_fifo_0_out_st_ready,                 //      tx_dma_fifo_0_out_st.ready
		output wire         tx_dma_fifo_0_out_st_startofpacket,         //                          .startofpacket
		output wire         tx_dma_fifo_0_out_st_valid,                 //                          .valid
		output wire         tx_dma_fifo_0_out_st_endofpacket,           //                          .endofpacket
		output wire [63:0]  tx_dma_fifo_0_out_st_data,                  //                          .data
		output wire [2:0]   tx_dma_fifo_0_out_st_empty,                 //                          .empty
		output wire [0:0]   tx_dma_fifo_0_out_st_error,                 //                          .error
		output wire         tx_dma_fifo_0_out_ts_req_valid,             //  tx_dma_fifo_0_out_ts_req.valid
		output wire [19:0]  tx_dma_fifo_0_out_ts_req_fingerprint,       //                          .fingerprint
		input  wire         ftile_clk_clk,                              //                 ftile_clk.clk
		output wire [36:0]  prefetcher_read_master_address,             //    prefetcher_read_master.address
		output wire         prefetcher_read_master_read,                //                          .read
		input  wire [127:0] prefetcher_read_master_readdata,            //                          .readdata
		input  wire         prefetcher_read_master_waitrequest,         //                          .waitrequest
		input  wire         prefetcher_read_master_readdatavalid,       //                          .readdatavalid
		output wire [2:0]   prefetcher_read_master_burstcount,          //                          .burstcount
		output wire [36:0]  prefetcher_write_master_address,            //   prefetcher_write_master.address
		output wire         prefetcher_write_master_write,              //                          .write
		output wire [15:0]  prefetcher_write_master_byteenable,         //                          .byteenable
		output wire [127:0] prefetcher_write_master_writedata,          //                          .writedata
		input  wire         prefetcher_write_master_waitrequest,        //                          .waitrequest
		input  wire [1:0]   prefetcher_write_master_response,           //                          .response
		input  wire         prefetcher_write_master_writeresponsevalid, //                          .writeresponsevalid
		output wire         irq_irq,                                    //                       irq.irq
		output wire [36:0]  read_master_address,                        //               read_master.address
		output wire         read_master_read,                           //                          .read
		output wire [15:0]  read_master_byteenable,                     //                          .byteenable
		input  wire [127:0] read_master_readdata,                       //                          .readdata
		input  wire         read_master_waitrequest,                    //                          .waitrequest
		input  wire         read_master_readdatavalid,                  //                          .readdatavalid
		output wire [4:0]   read_master_burstcount,                     //                          .burstcount
		input  wire         reset_reset_n                               //                     reset.reset_n
	);

	wire          tx_dma_prefetcher_descriptor_write_dispatcher_source_valid; // tx_dma_prefetcher:st_src_descr_valid -> tx_dma_dispatcher:snk_descriptor_valid
	wire  [255:0] tx_dma_prefetcher_descriptor_write_dispatcher_source_data;  // tx_dma_prefetcher:st_src_descr_data -> tx_dma_dispatcher:snk_descriptor_data
	wire          tx_dma_prefetcher_descriptor_write_dispatcher_source_ready; // tx_dma_dispatcher:snk_descriptor_ready -> tx_dma_prefetcher:st_src_descr_ready
	wire          tx_dma_dispatcher_read_command_source_valid;                // tx_dma_dispatcher:src_read_master_valid -> tx_dma_read_master:snk_command_valid
	wire  [255:0] tx_dma_dispatcher_read_command_source_data;                 // tx_dma_dispatcher:src_read_master_data -> tx_dma_read_master:snk_command_data
	wire          tx_dma_dispatcher_read_command_source_ready;                // tx_dma_read_master:snk_command_ready -> tx_dma_dispatcher:src_read_master_ready
	wire          tx_dma_read_master_response_source_valid;                   // tx_dma_read_master:src_response_valid -> tx_dma_dispatcher:snk_read_master_valid
	wire  [255:0] tx_dma_read_master_response_source_data;                    // tx_dma_read_master:src_response_data -> tx_dma_dispatcher:snk_read_master_data
	wire          tx_dma_read_master_response_source_ready;                   // tx_dma_dispatcher:snk_read_master_ready -> tx_dma_read_master:src_response_ready
	wire          tx_dma_dispatcher_response_source_valid;                    // tx_dma_dispatcher:src_response_valid -> tx_dma_fifo_0:in_ts_resp_valid
	wire  [255:0] tx_dma_dispatcher_response_source_data;                     // tx_dma_dispatcher:src_response_data -> tx_dma_fifo_0:in_ts_resp_data
	wire          tx_dma_dispatcher_response_source_ready;                    // tx_dma_fifo_0:in_ts_resp_ready -> tx_dma_dispatcher:src_response_ready
	wire          ts_chs_compl_0_out_st_valid;                                // ts_chs_compl_0:out_st_valid -> tx_dma_fifo_0:in_st_valid
	wire   [63:0] ts_chs_compl_0_out_st_data;                                 // ts_chs_compl_0:out_st_data -> tx_dma_fifo_0:in_st_data
	wire          ts_chs_compl_0_out_st_ready;                                // tx_dma_fifo_0:in_st_ready -> ts_chs_compl_0:out_st_ready
	wire          ts_chs_compl_0_out_st_startofpacket;                        // ts_chs_compl_0:out_st_sop -> tx_dma_fifo_0:in_st_sop
	wire          ts_chs_compl_0_out_st_endofpacket;                          // ts_chs_compl_0:out_st_eop -> tx_dma_fifo_0:in_st_eop
	wire          ts_chs_compl_0_out_st_error;                                // ts_chs_compl_0:out_st_error -> tx_dma_fifo_0:in_st_error
	wire    [2:0] ts_chs_compl_0_out_st_empty;                                // ts_chs_compl_0:out_st_empty -> tx_dma_fifo_0:in_st_empty
	wire          tx_dma_fifo_0_out_ts_resp_valid;                            // tx_dma_fifo_0:out_ts_resp_valid -> tx_dma_prefetcher:st_snk_valid
	wire  [255:0] tx_dma_fifo_0_out_ts_resp_data;                             // tx_dma_fifo_0:out_ts_resp_data -> tx_dma_prefetcher:st_snk_data
	wire          tx_dma_fifo_0_out_ts_resp_ready;                            // tx_dma_prefetcher:st_snk_ready -> tx_dma_fifo_0:out_ts_resp_ready
	wire          tx_dma_clock_out_clk_clk;                                   // tx_dma_clock:out_clk -> [avalon_st_adapter:in_clk_0_clk, mm_interconnect_0:tx_dma_clock_out_clk_clk, ts_chs_compl_0:i_ts_req_clk, tx_dma_csr:clk, tx_dma_dispatcher:clk, tx_dma_fifo_0:csr_clk, tx_dma_fifo_0:in_st_clk, tx_dma_fifo_0:ts_resp_clk, tx_dma_prefetcher:clk, tx_dma_read_master:clk, tx_dma_reset:clk]
	wire          tx_dma_ftile_clock_out_clk_clk;                             // tx_dma_ftile_clock:out_clk -> [rst_controller:clk, tx_dma_fifo_0:out_st_clk]
	wire    [0:0] ts_chs_compl_0_o_ts_valid;                                  // ts_chs_compl_0:o_ts_valid -> tx_dma_fifo_0:in_ts_valid
	wire   [95:0] ts_chs_compl_0_o_ts_data;                                   // ts_chs_compl_0:o_ts_data -> tx_dma_fifo_0:in_ts_data
	wire   [19:0] ts_chs_compl_0_o_ts_fingerprint;                            // ts_chs_compl_0:o_ts_fp -> tx_dma_fifo_0:in_ts_fp
	wire          tx_dma_reset_out_reset_reset;                               // tx_dma_reset:out_reset_n -> [avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:tx_dma_csr_reset_reset_bridge_in_reset_reset, mm_interconnect_0:tx_dma_dispatcher_clock_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0, ts_chs_compl_0:i_ts_req_rst, tx_dma_csr:reset, tx_dma_dispatcher:reset, tx_dma_fifo_0:csr_rst, tx_dma_fifo_0:in_st_rst, tx_dma_fifo_0:ts_resp_rst, tx_dma_prefetcher:reset, tx_dma_read_master:reset]
	wire          tx_dma_csr_m0_waitrequest;                                  // mm_interconnect_0:tx_dma_csr_m0_waitrequest -> tx_dma_csr:m0_waitrequest
	wire   [31:0] tx_dma_csr_m0_readdata;                                     // mm_interconnect_0:tx_dma_csr_m0_readdata -> tx_dma_csr:m0_readdata
	wire          tx_dma_csr_m0_debugaccess;                                  // tx_dma_csr:m0_debugaccess -> mm_interconnect_0:tx_dma_csr_m0_debugaccess
	wire    [5:0] tx_dma_csr_m0_address;                                      // tx_dma_csr:m0_address -> mm_interconnect_0:tx_dma_csr_m0_address
	wire          tx_dma_csr_m0_read;                                         // tx_dma_csr:m0_read -> mm_interconnect_0:tx_dma_csr_m0_read
	wire    [3:0] tx_dma_csr_m0_byteenable;                                   // tx_dma_csr:m0_byteenable -> mm_interconnect_0:tx_dma_csr_m0_byteenable
	wire          tx_dma_csr_m0_readdatavalid;                                // mm_interconnect_0:tx_dma_csr_m0_readdatavalid -> tx_dma_csr:m0_readdatavalid
	wire   [31:0] tx_dma_csr_m0_writedata;                                    // tx_dma_csr:m0_writedata -> mm_interconnect_0:tx_dma_csr_m0_writedata
	wire          tx_dma_csr_m0_write;                                        // tx_dma_csr:m0_write -> mm_interconnect_0:tx_dma_csr_m0_write
	wire    [0:0] tx_dma_csr_m0_burstcount;                                   // tx_dma_csr:m0_burstcount -> mm_interconnect_0:tx_dma_csr_m0_burstcount
	wire   [31:0] mm_interconnect_0_tx_dma_dispatcher_csr_readdata;           // tx_dma_dispatcher:csr_readdata -> mm_interconnect_0:tx_dma_dispatcher_CSR_readdata
	wire    [2:0] mm_interconnect_0_tx_dma_dispatcher_csr_address;            // mm_interconnect_0:tx_dma_dispatcher_CSR_address -> tx_dma_dispatcher:csr_address
	wire          mm_interconnect_0_tx_dma_dispatcher_csr_read;               // mm_interconnect_0:tx_dma_dispatcher_CSR_read -> tx_dma_dispatcher:csr_read
	wire    [3:0] mm_interconnect_0_tx_dma_dispatcher_csr_byteenable;         // mm_interconnect_0:tx_dma_dispatcher_CSR_byteenable -> tx_dma_dispatcher:csr_byteenable
	wire          mm_interconnect_0_tx_dma_dispatcher_csr_write;              // mm_interconnect_0:tx_dma_dispatcher_CSR_write -> tx_dma_dispatcher:csr_write
	wire   [31:0] mm_interconnect_0_tx_dma_dispatcher_csr_writedata;          // mm_interconnect_0:tx_dma_dispatcher_CSR_writedata -> tx_dma_dispatcher:csr_writedata
	wire   [31:0] mm_interconnect_0_tx_dma_prefetcher_csr_readdata;           // tx_dma_prefetcher:mm_csr_readdata -> mm_interconnect_0:tx_dma_prefetcher_Csr_readdata
	wire    [2:0] mm_interconnect_0_tx_dma_prefetcher_csr_address;            // mm_interconnect_0:tx_dma_prefetcher_Csr_address -> tx_dma_prefetcher:mm_csr_address
	wire          mm_interconnect_0_tx_dma_prefetcher_csr_read;               // mm_interconnect_0:tx_dma_prefetcher_Csr_read -> tx_dma_prefetcher:mm_csr_read
	wire          mm_interconnect_0_tx_dma_prefetcher_csr_write;              // mm_interconnect_0:tx_dma_prefetcher_Csr_write -> tx_dma_prefetcher:mm_csr_write
	wire   [31:0] mm_interconnect_0_tx_dma_prefetcher_csr_writedata;          // mm_interconnect_0:tx_dma_prefetcher_Csr_writedata -> tx_dma_prefetcher:mm_csr_writedata
	wire          tx_dma_read_master_data_source_valid;                       // tx_dma_read_master:src_valid -> avalon_st_adapter:in_0_valid
	wire  [127:0] tx_dma_read_master_data_source_data;                        // tx_dma_read_master:src_data -> avalon_st_adapter:in_0_data
	wire          tx_dma_read_master_data_source_ready;                       // avalon_st_adapter:in_0_ready -> tx_dma_read_master:src_ready
	wire          tx_dma_read_master_data_source_startofpacket;               // tx_dma_read_master:src_sop -> avalon_st_adapter:in_0_startofpacket
	wire          tx_dma_read_master_data_source_endofpacket;                 // tx_dma_read_master:src_eop -> avalon_st_adapter:in_0_endofpacket
	wire          tx_dma_read_master_data_source_error;                       // tx_dma_read_master:src_error -> avalon_st_adapter:in_0_error
	wire    [3:0] tx_dma_read_master_data_source_empty;                       // tx_dma_read_master:src_empty -> avalon_st_adapter:in_0_empty
	wire          avalon_st_adapter_out_0_valid;                              // avalon_st_adapter:out_0_valid -> ts_chs_compl_0:in_st_valid
	wire   [63:0] avalon_st_adapter_out_0_data;                               // avalon_st_adapter:out_0_data -> ts_chs_compl_0:in_st_data
	wire          avalon_st_adapter_out_0_ready;                              // ts_chs_compl_0:in_st_ready -> avalon_st_adapter:out_0_ready
	wire          avalon_st_adapter_out_0_startofpacket;                      // avalon_st_adapter:out_0_startofpacket -> ts_chs_compl_0:in_st_sop
	wire          avalon_st_adapter_out_0_endofpacket;                        // avalon_st_adapter:out_0_endofpacket -> ts_chs_compl_0:in_st_eop
	wire          avalon_st_adapter_out_0_error;                              // avalon_st_adapter:out_0_error -> ts_chs_compl_0:in_st_error
	wire    [2:0] avalon_st_adapter_out_0_empty;                              // avalon_st_adapter:out_0_empty -> ts_chs_compl_0:in_st_empty
	wire          rst_controller_reset_out_reset;                             // rst_controller:reset_out -> tx_dma_fifo_0:out_st_rst

	msgdma_ptp_subsys_8chs_ts_chs_compl_0 ts_chs_compl_0 (
		.i_ts_req_clk (tx_dma_clock_out_clk_clk),              //   input,   width = 1,   ts_req_clk.clk
		.i_ts_req_rst (~tx_dma_reset_out_reset_reset),         //   input,   width = 1, ts_req_reset.reset
		.i_clk_bus    (ts_chs_compl_0_clk_bus_in_clk),         //   input,   width = 1,   clk_bus_in.clk
		.i_rst_bus    (ts_chs_compl_0_rst_bus_in_reset),       //   input,   width = 1,   rst_bus_in.reset
		.in_st_ready  (avalon_st_adapter_out_0_ready),         //  output,   width = 1,        in_st.ready
		.in_st_sop    (avalon_st_adapter_out_0_startofpacket), //   input,   width = 1,             .startofpacket
		.in_st_valid  (avalon_st_adapter_out_0_valid),         //   input,   width = 1,             .valid
		.in_st_eop    (avalon_st_adapter_out_0_endofpacket),   //   input,   width = 1,             .endofpacket
		.in_st_data   (avalon_st_adapter_out_0_data),          //   input,  width = 64,             .data
		.in_st_empty  (avalon_st_adapter_out_0_empty),         //   input,   width = 3,             .empty
		.in_st_error  (avalon_st_adapter_out_0_error),         //   input,   width = 1,             .error
		.out_st_ready (ts_chs_compl_0_out_st_ready),           //   input,   width = 1,       out_st.ready
		.out_st_sop   (ts_chs_compl_0_out_st_startofpacket),   //  output,   width = 1,             .startofpacket
		.out_st_valid (ts_chs_compl_0_out_st_valid),           //  output,   width = 1,             .valid
		.out_st_eop   (ts_chs_compl_0_out_st_endofpacket),     //  output,   width = 1,             .endofpacket
		.out_st_data  (ts_chs_compl_0_out_st_data),            //  output,  width = 64,             .data
		.out_st_empty (ts_chs_compl_0_out_st_empty),           //  output,   width = 3,             .empty
		.out_st_error (ts_chs_compl_0_out_st_error),           //  output,   width = 1,             .error
		.i_ts_valid   (ts_chs_compl_0_i_ts_valid),             //   input,   width = 1,         i_ts.valid
		.i_ts_fp      (ts_chs_compl_0_i_ts_fingerprint),       //   input,  width = 20,             .fingerprint
		.i_ts_data    (ts_chs_compl_0_i_ts_data),              //   input,  width = 96,             .data
		.o_ts_valid   (ts_chs_compl_0_o_ts_valid),             //  output,   width = 1,         o_ts.valid
		.o_ts_fp      (ts_chs_compl_0_o_ts_fingerprint),       //  output,  width = 20,             .fingerprint
		.o_ts_data    (ts_chs_compl_0_o_ts_data)               //  output,  width = 96,             .data
	);

	tx_dma_clock tx_dma_clock (
		.in_clk  (dma_clk_clk),              //   input,  width = 1,  in_clk.clk
		.out_clk (tx_dma_clock_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	tx_dma_csr tx_dma_csr (
		.clk              (tx_dma_clock_out_clk_clk),      //   input,   width = 1,   clk.clk
		.reset            (~tx_dma_reset_out_reset_reset), //   input,   width = 1, reset.reset
		.s0_waitrequest   (csr_waitrequest),               //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (csr_readdata),                  //  output,  width = 32,      .readdata
		.s0_readdatavalid (csr_readdatavalid),             //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (csr_burstcount),                //   input,   width = 1,      .burstcount
		.s0_writedata     (csr_writedata),                 //   input,  width = 32,      .writedata
		.s0_address       (csr_address),                   //   input,   width = 6,      .address
		.s0_write         (csr_write),                     //   input,   width = 1,      .write
		.s0_read          (csr_read),                      //   input,   width = 1,      .read
		.s0_byteenable    (csr_byteenable),                //   input,   width = 4,      .byteenable
		.s0_debugaccess   (csr_debugaccess),               //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (tx_dma_csr_m0_waitrequest),     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (tx_dma_csr_m0_readdata),        //   input,  width = 32,      .readdata
		.m0_readdatavalid (tx_dma_csr_m0_readdatavalid),   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (tx_dma_csr_m0_burstcount),      //  output,   width = 1,      .burstcount
		.m0_writedata     (tx_dma_csr_m0_writedata),       //  output,  width = 32,      .writedata
		.m0_address       (tx_dma_csr_m0_address),         //  output,   width = 6,      .address
		.m0_write         (tx_dma_csr_m0_write),           //  output,   width = 1,      .write
		.m0_read          (tx_dma_csr_m0_read),            //  output,   width = 1,      .read
		.m0_byteenable    (tx_dma_csr_m0_byteenable),      //  output,   width = 4,      .byteenable
		.m0_debugaccess   (tx_dma_csr_m0_debugaccess)      //  output,   width = 1,      .debugaccess
	);

	tx_dma_dispatcher tx_dma_dispatcher (
		.clk                   (tx_dma_clock_out_clk_clk),                                   //   input,    width = 1,               clock.clk
		.reset                 (~tx_dma_reset_out_reset_reset),                              //   input,    width = 1,         clock_reset.reset
		.csr_writedata         (mm_interconnect_0_tx_dma_dispatcher_csr_writedata),          //   input,   width = 32,                 CSR.writedata
		.csr_write             (mm_interconnect_0_tx_dma_dispatcher_csr_write),              //   input,    width = 1,                    .write
		.csr_byteenable        (mm_interconnect_0_tx_dma_dispatcher_csr_byteenable),         //   input,    width = 4,                    .byteenable
		.csr_readdata          (mm_interconnect_0_tx_dma_dispatcher_csr_readdata),           //  output,   width = 32,                    .readdata
		.csr_read              (mm_interconnect_0_tx_dma_dispatcher_csr_read),               //   input,    width = 1,                    .read
		.csr_address           (mm_interconnect_0_tx_dma_dispatcher_csr_address),            //   input,    width = 3,                    .address
		.src_response_data     (tx_dma_dispatcher_response_source_data),                     //  output,  width = 256,     Response_Source.data
		.src_response_valid    (tx_dma_dispatcher_response_source_valid),                    //  output,    width = 1,                    .valid
		.src_response_ready    (tx_dma_dispatcher_response_source_ready),                    //   input,    width = 1,                    .ready
		.snk_descriptor_data   (tx_dma_prefetcher_descriptor_write_dispatcher_source_data),  //   input,  width = 256,     Descriptor_Sink.data
		.snk_descriptor_valid  (tx_dma_prefetcher_descriptor_write_dispatcher_source_valid), //   input,    width = 1,                    .valid
		.snk_descriptor_ready  (tx_dma_prefetcher_descriptor_write_dispatcher_source_ready), //  output,    width = 1,                    .ready
		.src_read_master_data  (tx_dma_dispatcher_read_command_source_data),                 //  output,  width = 256, Read_Command_Source.data
		.src_read_master_valid (tx_dma_dispatcher_read_command_source_valid),                //  output,    width = 1,                    .valid
		.src_read_master_ready (tx_dma_dispatcher_read_command_source_ready),                //   input,    width = 1,                    .ready
		.snk_read_master_data  (tx_dma_read_master_response_source_data),                    //   input,  width = 256,  Read_Response_Sink.data
		.snk_read_master_valid (tx_dma_read_master_response_source_valid),                   //   input,    width = 1,                    .valid
		.snk_read_master_ready (tx_dma_read_master_response_source_ready)                    //  output,    width = 1,                    .ready
	);

	tx_dma_fifo_0 #(
		.DEVICE                ("s10"),
		.USE_RX_READY          (1),
		.MEMORY_CAPACITY_WORDS (1024),
		.AVST_DATA_WIDTH       (64),
		.AVST_ERROR_WIDTH      (1),
		.TS_FIFOS_ADDR_WIDTH   (9),
		.TS_WIDTH              (96),
		.TS_RESP_WIDTH         (256),
		.TS_FP_WIDTH           (20),
		.AVST_EMPTY_WIDTH      (3),
		.DEBUG_EN              (1)
	) tx_dma_fifo_0 (
		.in_st_clk              (tx_dma_clock_out_clk_clk),                //   input,    width = 1,   in_st_clk.clk
		.in_st_rst              (~tx_dma_reset_out_reset_reset),           //   input,    width = 1,   in_st_rst.reset
		.out_st_clk             (tx_dma_ftile_clock_out_clk_clk),          //   input,    width = 1,  out_st_clk.clk
		.out_st_rst             (rst_controller_reset_out_reset),          //   input,    width = 1,  out_st_rst.reset
		.ts_resp_clk            (tx_dma_clock_out_clk_clk),                //   input,    width = 1, ts_resp_clk.clk
		.ts_resp_rst            (~tx_dma_reset_out_reset_reset),           //   input,    width = 1, ts_resp_rst.reset
		.csr_clk                (tx_dma_clock_out_clk_clk),                //   input,    width = 1,     csr_clk.clk
		.csr_rst                (~tx_dma_reset_out_reset_reset),           //   input,    width = 1,     csr_rst.reset
		.in_st_ready            (ts_chs_compl_0_out_st_ready),             //  output,    width = 1,       in_st.ready
		.in_st_sop              (ts_chs_compl_0_out_st_startofpacket),     //   input,    width = 1,            .startofpacket
		.in_st_valid            (ts_chs_compl_0_out_st_valid),             //   input,    width = 1,            .valid
		.in_st_eop              (ts_chs_compl_0_out_st_endofpacket),       //   input,    width = 1,            .endofpacket
		.in_st_data             (ts_chs_compl_0_out_st_data),              //   input,   width = 64,            .data
		.in_st_empty            (ts_chs_compl_0_out_st_empty),             //   input,    width = 3,            .empty
		.in_st_error            (ts_chs_compl_0_out_st_error),             //   input,    width = 1,            .error
		.out_st_ready           (tx_dma_fifo_0_out_st_ready),              //   input,    width = 1,      out_st.ready
		.out_st_sop             (tx_dma_fifo_0_out_st_startofpacket),      //  output,    width = 1,            .startofpacket
		.out_st_valid           (tx_dma_fifo_0_out_st_valid),              //  output,    width = 1,            .valid
		.out_st_eop             (tx_dma_fifo_0_out_st_endofpacket),        //  output,    width = 1,            .endofpacket
		.out_st_data            (tx_dma_fifo_0_out_st_data),               //  output,   width = 64,            .data
		.out_st_empty           (tx_dma_fifo_0_out_st_empty),              //  output,    width = 3,            .empty
		.out_st_error           (tx_dma_fifo_0_out_st_error),              //  output,    width = 1,            .error
		.in_ts_resp_ready       (tx_dma_dispatcher_response_source_ready), //  output,    width = 1,  in_ts_resp.ready
		.in_ts_resp_valid       (tx_dma_dispatcher_response_source_valid), //   input,    width = 1,            .valid
		.in_ts_resp_data        (tx_dma_dispatcher_response_source_data),  //   input,  width = 256,            .data
		.out_ts_resp_ready      (tx_dma_fifo_0_out_ts_resp_ready),         //   input,    width = 1, out_ts_resp.ready
		.out_ts_resp_valid      (tx_dma_fifo_0_out_ts_resp_valid),         //  output,    width = 1,            .valid
		.out_ts_resp_data       (tx_dma_fifo_0_out_ts_resp_data),          //  output,  width = 256,            .data
		.out_ts_req_valid       (tx_dma_fifo_0_out_ts_req_valid),          //  output,    width = 1,  out_ts_req.valid
		.out_ts_req_fingerprint (tx_dma_fifo_0_out_ts_req_fingerprint),    //  output,   width = 20,            .fingerprint
		.in_ts_valid            (ts_chs_compl_0_o_ts_valid),               //   input,    width = 1,       in_ts.valid
		.in_ts_fp               (ts_chs_compl_0_o_ts_fingerprint),         //   input,   width = 20,            .fingerprint
		.in_ts_data             (ts_chs_compl_0_o_ts_data)                 //   input,   width = 96,            .data
	);

	tx_dma_ftile_clock tx_dma_ftile_clock (
		.in_clk  (ftile_clk_clk),                  //   input,  width = 1,  in_clk.clk
		.out_clk (tx_dma_ftile_clock_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	tx_dma_prefetcher tx_dma_prefetcher (
		.clk                         (tx_dma_clock_out_clk_clk),                                   //   input,    width = 1,                              Clock.clk
		.reset                       (~tx_dma_reset_out_reset_reset),                              //   input,    width = 1,                        Clock_reset.reset
		.mm_read_address             (prefetcher_read_master_address),                             //  output,   width = 37,             Descriptor_Read_Master.address
		.mm_read_read                (prefetcher_read_master_read),                                //  output,    width = 1,                                   .read
		.mm_read_readdata            (prefetcher_read_master_readdata),                            //   input,  width = 128,                                   .readdata
		.mm_read_waitrequest         (prefetcher_read_master_waitrequest),                         //   input,    width = 1,                                   .waitrequest
		.mm_read_readdatavalid       (prefetcher_read_master_readdatavalid),                       //   input,    width = 1,                                   .readdatavalid
		.mm_read_burstcount          (prefetcher_read_master_burstcount),                          //  output,    width = 3,                                   .burstcount
		.mm_write_address            (prefetcher_write_master_address),                            //  output,   width = 37,            Descriptor_Write_Master.address
		.mm_write_write              (prefetcher_write_master_write),                              //  output,    width = 1,                                   .write
		.mm_write_byteenable         (prefetcher_write_master_byteenable),                         //  output,   width = 16,                                   .byteenable
		.mm_write_writedata          (prefetcher_write_master_writedata),                          //  output,  width = 128,                                   .writedata
		.mm_write_waitrequest        (prefetcher_write_master_waitrequest),                        //   input,    width = 1,                                   .waitrequest
		.mm_write_response           (prefetcher_write_master_response),                           //   input,    width = 2,                                   .response
		.mm_write_writeresponsevalid (prefetcher_write_master_writeresponsevalid),                 //   input,    width = 1,                                   .writeresponsevalid
		.st_src_descr_data           (tx_dma_prefetcher_descriptor_write_dispatcher_source_data),  //  output,  width = 256, Descriptor_Write_Dispatcher_Source.data
		.st_src_descr_valid          (tx_dma_prefetcher_descriptor_write_dispatcher_source_valid), //  output,    width = 1,                                   .valid
		.st_src_descr_ready          (tx_dma_prefetcher_descriptor_write_dispatcher_source_ready), //   input,    width = 1,                                   .ready
		.st_snk_data                 (tx_dma_fifo_0_out_ts_resp_data),                             //   input,  width = 256,                      Response_Sink.data
		.st_snk_valid                (tx_dma_fifo_0_out_ts_resp_valid),                            //   input,    width = 1,                                   .valid
		.st_snk_ready                (tx_dma_fifo_0_out_ts_resp_ready),                            //  output,    width = 1,                                   .ready
		.mm_csr_address              (mm_interconnect_0_tx_dma_prefetcher_csr_address),            //   input,    width = 3,                                Csr.address
		.mm_csr_read                 (mm_interconnect_0_tx_dma_prefetcher_csr_read),               //   input,    width = 1,                                   .read
		.mm_csr_write                (mm_interconnect_0_tx_dma_prefetcher_csr_write),              //   input,    width = 1,                                   .write
		.mm_csr_writedata            (mm_interconnect_0_tx_dma_prefetcher_csr_writedata),          //   input,   width = 32,                                   .writedata
		.mm_csr_readdata             (mm_interconnect_0_tx_dma_prefetcher_csr_readdata),           //  output,   width = 32,                                   .readdata
		.csr_irq                     (irq_irq)                                                     //  output,    width = 1,                            Csr_Irq.irq
	);

	tx_dma_read_master tx_dma_read_master (
		.clk                  (tx_dma_clock_out_clk_clk),                     //   input,    width = 1,            Clock.clk
		.reset                (~tx_dma_reset_out_reset_reset),                //   input,    width = 1,      Clock_reset.reset
		.master_address       (read_master_address),                          //  output,   width = 37, Data_Read_Master.address
		.master_read          (read_master_read),                             //  output,    width = 1,                 .read
		.master_byteenable    (read_master_byteenable),                       //  output,   width = 16,                 .byteenable
		.master_readdata      (read_master_readdata),                         //   input,  width = 128,                 .readdata
		.master_waitrequest   (read_master_waitrequest),                      //   input,    width = 1,                 .waitrequest
		.master_readdatavalid (read_master_readdatavalid),                    //   input,    width = 1,                 .readdatavalid
		.master_burstcount    (read_master_burstcount),                       //  output,    width = 5,                 .burstcount
		.src_data             (tx_dma_read_master_data_source_data),          //  output,  width = 128,      Data_Source.data
		.src_valid            (tx_dma_read_master_data_source_valid),         //  output,    width = 1,                 .valid
		.src_ready            (tx_dma_read_master_data_source_ready),         //   input,    width = 1,                 .ready
		.src_sop              (tx_dma_read_master_data_source_startofpacket), //  output,    width = 1,                 .startofpacket
		.src_eop              (tx_dma_read_master_data_source_endofpacket),   //  output,    width = 1,                 .endofpacket
		.src_empty            (tx_dma_read_master_data_source_empty),         //  output,    width = 4,                 .empty
		.src_error            (tx_dma_read_master_data_source_error),         //  output,    width = 1,                 .error
		.snk_command_data     (tx_dma_dispatcher_read_command_source_data),   //   input,  width = 256,     Command_Sink.data
		.snk_command_valid    (tx_dma_dispatcher_read_command_source_valid),  //   input,    width = 1,                 .valid
		.snk_command_ready    (tx_dma_dispatcher_read_command_source_ready),  //  output,    width = 1,                 .ready
		.src_response_data    (tx_dma_read_master_response_source_data),      //  output,  width = 256,  Response_Source.data
		.src_response_valid   (tx_dma_read_master_response_source_valid),     //  output,    width = 1,                 .valid
		.src_response_ready   (tx_dma_read_master_response_source_ready)      //   input,    width = 1,                 .ready
	);

	tx_dma_reset tx_dma_reset (
		.clk         (tx_dma_clock_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_reset_n),                //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (tx_dma_reset_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	subsys_ftile_25gbe_tx_dma_altera_mm_interconnect_1920_4olduea mm_interconnect_0 (
		.tx_dma_csr_m0_address                                     (tx_dma_csr_m0_address),                              //   input,   width = 6,                                       tx_dma_csr_m0.address
		.tx_dma_csr_m0_waitrequest                                 (tx_dma_csr_m0_waitrequest),                          //  output,   width = 1,                                                    .waitrequest
		.tx_dma_csr_m0_burstcount                                  (tx_dma_csr_m0_burstcount),                           //   input,   width = 1,                                                    .burstcount
		.tx_dma_csr_m0_byteenable                                  (tx_dma_csr_m0_byteenable),                           //   input,   width = 4,                                                    .byteenable
		.tx_dma_csr_m0_read                                        (tx_dma_csr_m0_read),                                 //   input,   width = 1,                                                    .read
		.tx_dma_csr_m0_readdata                                    (tx_dma_csr_m0_readdata),                             //  output,  width = 32,                                                    .readdata
		.tx_dma_csr_m0_readdatavalid                               (tx_dma_csr_m0_readdatavalid),                        //  output,   width = 1,                                                    .readdatavalid
		.tx_dma_csr_m0_write                                       (tx_dma_csr_m0_write),                                //   input,   width = 1,                                                    .write
		.tx_dma_csr_m0_writedata                                   (tx_dma_csr_m0_writedata),                            //   input,  width = 32,                                                    .writedata
		.tx_dma_csr_m0_debugaccess                                 (tx_dma_csr_m0_debugaccess),                          //   input,   width = 1,                                                    .debugaccess
		.tx_dma_dispatcher_CSR_address                             (mm_interconnect_0_tx_dma_dispatcher_csr_address),    //  output,   width = 3,                               tx_dma_dispatcher_CSR.address
		.tx_dma_dispatcher_CSR_write                               (mm_interconnect_0_tx_dma_dispatcher_csr_write),      //  output,   width = 1,                                                    .write
		.tx_dma_dispatcher_CSR_read                                (mm_interconnect_0_tx_dma_dispatcher_csr_read),       //  output,   width = 1,                                                    .read
		.tx_dma_dispatcher_CSR_readdata                            (mm_interconnect_0_tx_dma_dispatcher_csr_readdata),   //   input,  width = 32,                                                    .readdata
		.tx_dma_dispatcher_CSR_writedata                           (mm_interconnect_0_tx_dma_dispatcher_csr_writedata),  //  output,  width = 32,                                                    .writedata
		.tx_dma_dispatcher_CSR_byteenable                          (mm_interconnect_0_tx_dma_dispatcher_csr_byteenable), //  output,   width = 4,                                                    .byteenable
		.tx_dma_prefetcher_Csr_address                             (mm_interconnect_0_tx_dma_prefetcher_csr_address),    //  output,   width = 3,                               tx_dma_prefetcher_Csr.address
		.tx_dma_prefetcher_Csr_write                               (mm_interconnect_0_tx_dma_prefetcher_csr_write),      //  output,   width = 1,                                                    .write
		.tx_dma_prefetcher_Csr_read                                (mm_interconnect_0_tx_dma_prefetcher_csr_read),       //  output,   width = 1,                                                    .read
		.tx_dma_prefetcher_Csr_readdata                            (mm_interconnect_0_tx_dma_prefetcher_csr_readdata),   //   input,  width = 32,                                                    .readdata
		.tx_dma_prefetcher_Csr_writedata                           (mm_interconnect_0_tx_dma_prefetcher_csr_writedata),  //  output,  width = 32,                                                    .writedata
		.tx_dma_csr_reset_reset_bridge_in_reset_reset              (~tx_dma_reset_out_reset_reset),                      //   input,   width = 1,              tx_dma_csr_reset_reset_bridge_in_reset.reset
		.tx_dma_dispatcher_clock_reset_reset_bridge_in_reset_reset (~tx_dma_reset_out_reset_reset),                      //   input,   width = 1, tx_dma_dispatcher_clock_reset_reset_bridge_in_reset.reset
		.tx_dma_clock_out_clk_clk                                  (tx_dma_clock_out_clk_clk)                            //   input,   width = 1,                                tx_dma_clock_out_clk.clk
	);

	subsys_ftile_25gbe_tx_dma_altera_avalon_st_adapter_1920_whdx2tq #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (128),
		.inChannelWidth  (0),
		.inErrorWidth    (1),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (64),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (tx_dma_clock_out_clk_clk),                     //   input,    width = 1, in_clk_0.clk
		.in_rst_0_reset      (~tx_dma_reset_out_reset_reset),                //   input,    width = 1, in_rst_0.reset
		.in_0_data           (tx_dma_read_master_data_source_data),          //   input,  width = 128,     in_0.data
		.in_0_valid          (tx_dma_read_master_data_source_valid),         //   input,    width = 1,         .valid
		.in_0_ready          (tx_dma_read_master_data_source_ready),         //  output,    width = 1,         .ready
		.in_0_startofpacket  (tx_dma_read_master_data_source_startofpacket), //   input,    width = 1,         .startofpacket
		.in_0_endofpacket    (tx_dma_read_master_data_source_endofpacket),   //   input,    width = 1,         .endofpacket
		.in_0_empty          (tx_dma_read_master_data_source_empty),         //   input,    width = 4,         .empty
		.in_0_error          (tx_dma_read_master_data_source_error),         //   input,    width = 1,         .error
		.out_0_data          (avalon_st_adapter_out_0_data),                 //  output,   width = 64,    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                //  output,    width = 1,         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                //   input,    width = 1,         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),        //  output,    width = 1,         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),          //  output,    width = 1,         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),                //  output,    width = 3,         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)                 //  output,    width = 1,         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~tx_dma_reset_out_reset_reset),  //   input,  width = 1, reset_in0.reset
		.clk            (tx_dma_ftile_clock_out_clk_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

endmodule
