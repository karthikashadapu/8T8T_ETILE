// dma_subsystem.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module dma_subsystem (
		output wire         acp_bridge_in_clk_clk,                                                        //                                                acp_bridge_in_clk.clk
		input  wire         dma_clk_100_in_clk_clk,                                                       //                                               dma_clk_100_in_clk.clk
		output wire         dma_clk_out_bridge_0_out_clk_clk,                                             //                                     dma_clk_out_bridge_0_out_clk.clk
		input  wire         dma_rst_100_in_reset_reset,                                                   //                                             dma_rst_100_in_reset.reset
		input  wire         dma_ss_master_m0_waitrequest,                                                 //                                                 dma_ss_master_m0.waitrequest
		input  wire [511:0] dma_ss_master_m0_readdata,                                                    //                                                                 .readdata
		input  wire         dma_ss_master_m0_readdatavalid,                                               //                                                                 .readdatavalid
		input  wire [1:0]   dma_ss_master_m0_response,                                                    //                                                                 .response
		output wire [4:0]   dma_ss_master_m0_burstcount,                                                  //                                                                 .burstcount
		output wire [511:0] dma_ss_master_m0_writedata,                                                   //                                                                 .writedata
		output wire [36:0]  dma_ss_master_m0_address,                                                     //                                                                 .address
		output wire         dma_ss_master_m0_write,                                                       //                                                                 .write
		output wire         dma_ss_master_m0_read,                                                        //                                                                 .read
		output wire [63:0]  dma_ss_master_m0_byteenable,                                                  //                                                                 .byteenable
		output wire         dma_ss_master_m0_debugaccess,                                                 //                                                                 .debugaccess
		input  wire         dma_ss_master_m0_writeresponsevalid,                                          //                                                                 .writeresponsevalid
		input  wire [29:0]  ext_hps_m_master_windowed_slave_address,                                      //                                  ext_hps_m_master_windowed_slave.address
		input  wire         ext_hps_m_master_windowed_slave_read,                                         //                                                                 .read
		output wire [31:0]  ext_hps_m_master_windowed_slave_readdata,                                     //                                                                 .readdata
		input  wire         ext_hps_m_master_windowed_slave_write,                                        //                                                                 .write
		input  wire [31:0]  ext_hps_m_master_windowed_slave_writedata,                                    //                                                                 .writedata
		output wire         ext_hps_m_master_windowed_slave_readdatavalid,                                //                                                                 .readdatavalid
		output wire         ext_hps_m_master_windowed_slave_waitrequest,                                  //                                                                 .waitrequest
		input  wire [3:0]   ext_hps_m_master_windowed_slave_byteenable,                                   //                                                                 .byteenable
		input  wire [0:0]   ext_hps_m_master_windowed_slave_burstcount,                                   //                                                                 .burstcount
		output wire [36:0]  ext_hps_m_master_expanded_master_address,                                     //                                 ext_hps_m_master_expanded_master.address
		output wire         ext_hps_m_master_expanded_master_read,                                        //                                                                 .read
		input  wire         ext_hps_m_master_expanded_master_waitrequest,                                 //                                                                 .waitrequest
		input  wire [31:0]  ext_hps_m_master_expanded_master_readdata,                                    //                                                                 .readdata
		output wire         ext_hps_m_master_expanded_master_write,                                       //                                                                 .write
		output wire [31:0]  ext_hps_m_master_expanded_master_writedata,                                   //                                                                 .writedata
		input  wire         ext_hps_m_master_expanded_master_readdatavalid,                               //                                                                 .readdatavalid
		output wire [3:0]   ext_hps_m_master_expanded_master_byteenable,                                  //                                                                 .byteenable
		output wire [0:0]   ext_hps_m_master_expanded_master_burstcount,                                  //                                                                 .burstcount
		input  wire         oclk_pll_port8_in_clk_clk,                                                    //                                            oclk_pll_port8_in_clk.clk
		input  wire         rx_dma_reset_bridge_0_in_reset_reset_n,                                       //                                   rx_dma_reset_bridge_0_in_reset.reset_n
		input  wire         rx_dma_reset_bridge_1_in_reset_reset_n,                                       //                                   rx_dma_reset_bridge_1_in_reset.reset_n
		output wire         subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset_reset_n,                    //                subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset.reset_n
		input  wire         ninit_done_reset,                                                             //                                                       ninit_done.reset
		output wire         dma_subsys_port8_csr_waitrequest,                                             //                                             dma_subsys_port8_csr.waitrequest
		output wire [31:0]  dma_subsys_port8_csr_readdata,                                                //                                                                 .readdata
		output wire         dma_subsys_port8_csr_readdatavalid,                                           //                                                                 .readdatavalid
		input  wire [0:0]   dma_subsys_port8_csr_burstcount,                                              //                                                                 .burstcount
		input  wire [31:0]  dma_subsys_port8_csr_writedata,                                               //                                                                 .writedata
		input  wire [7:0]   dma_subsys_port8_csr_address,                                                 //                                                                 .address
		input  wire         dma_subsys_port8_csr_write,                                                   //                                                                 .write
		input  wire         dma_subsys_port8_csr_read,                                                    //                                                                 .read
		input  wire [3:0]   dma_subsys_port8_csr_byteenable,                                              //                                                                 .byteenable
		input  wire         dma_subsys_port8_csr_debugaccess,                                             //                                                                 .debugaccess
		input  wire         dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_startofpacket,                  //                    dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin.startofpacket
		input  wire         dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_valid,                          //                                                                 .valid
		input  wire         dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_endofpacket,                    //                                                                 .endofpacket
		input  wire [63:0]  dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_data,                           //                                                                 .data
		input  wire [2:0]   dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_empty,                          //                                                                 .empty
		input  wire [5:0]   dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_error,                          //                                                                 .error
		input  wire         dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_valid,            //      dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts.valid
		input  wire [95:0]  dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_data,             //                                                                 .data
		output wire         dma_subsys_port8_rx_dma_ch1_irq_irq,                                          //                                  dma_subsys_port8_rx_dma_ch1_irq.irq
		input  wire [0:0]   dma_subsys_port8_ts_chs_compl_0_clk_bus_in_clk,                               //                       dma_subsys_port8_ts_chs_compl_0_clk_bus_in.clk
		input  wire [0:0]   dma_subsys_port8_ts_chs_compl_0_rst_bus_in_reset,                             //                       dma_subsys_port8_ts_chs_compl_0_rst_bus_in.reset
		input  wire [0:0]   dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_valid,            //      dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts.valid
		input  wire [19:0]  dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_fingerprint,      //                                                                 .fingerprint
		input  wire [95:0]  dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_data,             //                                                                 .data
		input  wire         dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready,           //     dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st.ready
		output wire         dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket,   //                                                                 .startofpacket
		output wire         dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid,           //                                                                 .valid
		output wire         dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket,     //                                                                 .endofpacket
		output wire [63:0]  dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data,            //                                                                 .data
		output wire [2:0]   dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty,           //                                                                 .empty
		output wire [0:0]   dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error,           //                                                                 .error
		output wire         dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_valid,       // dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req.valid
		output wire [19:0]  dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_fingerprint, //                                                                 .fingerprint
		output wire         dma_subsys_port8_tx_dma_ch1_irq_irq                                           //                                  dma_subsys_port8_tx_dma_ch1_irq.irq
	);

	wire          dma_clk_100_out_clk_clk;                                                // dma_clk_100:out_clk -> [dma_rst_100:clk, dma_subsys_port8:clk_clk, ext_hps_m_master:clk, rst_controller_003:clk, rx_dma_reset_bridge_0:clk, rx_dma_reset_bridge_1:clk]
	wire          oclk_pll_port8_out_clk_clk;                                             // oclk_pll_port8:out_clk -> [dma_subsys_port8:subsys_ftile_25gbe_1588_o_pll_clk_in_clk_clk, iopll_clk_avst_div2:refclk]
	wire          iopll_clk_avst_div2_outclk0_clk;                                        // iopll_clk_avst_div2:outclk_0 -> [acp_bridge_in_clk:in_clk, dma_clk_out_bridge_0:in_clk, dma_ss_master:clk, dma_subsys_port8:subsys_ftile_25gbe_1588_dmaclkout_in_clk_clk, mm_interconnect_0:iopll_clk_avst_div2_outclk0_clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk, rst_controller_004:clk, subsys_ftile_25gbe_1588_dmaclkout_reset:clk]
	wire          subsys_ftile_25gbe_1588_ninitdone_reset_out_reset_reset;                // subsys_ftile_25gbe_1588_ninitdone_reset:out_reset -> [iopll_clk_avst_div2:rst, rst_controller_001:reset_in0]
	wire          dma_rst_100_out_reset_reset;                                            // dma_rst_100:out_reset -> [ext_hps_m_master:reset, rst_controller:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0]
	wire  [127:0] dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdata;            // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdata -> dma_subsys_port8:rx_dma_ch1_prefetcher_read_master_readdata
	wire          dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_waitrequest;         // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_waitrequest -> dma_subsys_port8:rx_dma_ch1_prefetcher_read_master_waitrequest
	wire   [36:0] dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_address;             // dma_subsys_port8:rx_dma_ch1_prefetcher_read_master_address -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_address
	wire          dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_read;                // dma_subsys_port8:rx_dma_ch1_prefetcher_read_master_read -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_read
	wire          dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdatavalid;       // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdatavalid -> dma_subsys_port8:rx_dma_ch1_prefetcher_read_master_readdatavalid
	wire    [2:0] dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_burstcount;          // dma_subsys_port8:rx_dma_ch1_prefetcher_read_master_burstcount -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_burstcount
	wire          dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_waitrequest;        // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_waitrequest -> dma_subsys_port8:rx_dma_ch1_prefetcher_write_master_waitrequest
	wire   [36:0] dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_address;            // dma_subsys_port8:rx_dma_ch1_prefetcher_write_master_address -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_address
	wire   [15:0] dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_byteenable;         // dma_subsys_port8:rx_dma_ch1_prefetcher_write_master_byteenable -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_byteenable
	wire    [1:0] dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_response;           // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_response -> dma_subsys_port8:rx_dma_ch1_prefetcher_write_master_response
	wire          dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_write;              // dma_subsys_port8:rx_dma_ch1_prefetcher_write_master_write -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_write
	wire  [127:0] dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writedata;          // dma_subsys_port8:rx_dma_ch1_prefetcher_write_master_writedata -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writedata
	wire          dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writeresponsevalid; // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writeresponsevalid -> dma_subsys_port8:rx_dma_ch1_prefetcher_write_master_writeresponsevalid
	wire          dma_subsys_port8_rx_dma_ch1_write_master_waitrequest;                   // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_write_master_waitrequest -> dma_subsys_port8:rx_dma_ch1_write_master_waitrequest
	wire   [36:0] dma_subsys_port8_rx_dma_ch1_write_master_address;                       // dma_subsys_port8:rx_dma_ch1_write_master_address -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_write_master_address
	wire   [15:0] dma_subsys_port8_rx_dma_ch1_write_master_byteenable;                    // dma_subsys_port8:rx_dma_ch1_write_master_byteenable -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_write_master_byteenable
	wire    [1:0] dma_subsys_port8_rx_dma_ch1_write_master_response;                      // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_write_master_response -> dma_subsys_port8:rx_dma_ch1_write_master_response
	wire          dma_subsys_port8_rx_dma_ch1_write_master_write;                         // dma_subsys_port8:rx_dma_ch1_write_master_write -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_write_master_write
	wire  [127:0] dma_subsys_port8_rx_dma_ch1_write_master_writedata;                     // dma_subsys_port8:rx_dma_ch1_write_master_writedata -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_write_master_writedata
	wire          dma_subsys_port8_rx_dma_ch1_write_master_writeresponsevalid;            // mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_write_master_writeresponsevalid -> dma_subsys_port8:rx_dma_ch1_write_master_writeresponsevalid
	wire    [4:0] dma_subsys_port8_rx_dma_ch1_write_master_burstcount;                    // dma_subsys_port8:rx_dma_ch1_write_master_burstcount -> mm_interconnect_0:dma_subsys_port8_rx_dma_ch1_write_master_burstcount
	wire  [127:0] dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdata;            // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdata -> dma_subsys_port8:tx_dma_ch1_prefetcher_read_master_readdata
	wire          dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_waitrequest;         // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_waitrequest -> dma_subsys_port8:tx_dma_ch1_prefetcher_read_master_waitrequest
	wire   [36:0] dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_address;             // dma_subsys_port8:tx_dma_ch1_prefetcher_read_master_address -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_address
	wire          dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_read;                // dma_subsys_port8:tx_dma_ch1_prefetcher_read_master_read -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_read
	wire          dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdatavalid;       // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdatavalid -> dma_subsys_port8:tx_dma_ch1_prefetcher_read_master_readdatavalid
	wire    [2:0] dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_burstcount;          // dma_subsys_port8:tx_dma_ch1_prefetcher_read_master_burstcount -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_burstcount
	wire          dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_waitrequest;        // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_waitrequest -> dma_subsys_port8:tx_dma_ch1_prefetcher_write_master_waitrequest
	wire   [36:0] dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_address;            // dma_subsys_port8:tx_dma_ch1_prefetcher_write_master_address -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_address
	wire   [15:0] dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_byteenable;         // dma_subsys_port8:tx_dma_ch1_prefetcher_write_master_byteenable -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_byteenable
	wire    [1:0] dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_response;           // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_response -> dma_subsys_port8:tx_dma_ch1_prefetcher_write_master_response
	wire          dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_write;              // dma_subsys_port8:tx_dma_ch1_prefetcher_write_master_write -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_write
	wire  [127:0] dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writedata;          // dma_subsys_port8:tx_dma_ch1_prefetcher_write_master_writedata -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writedata
	wire          dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writeresponsevalid; // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writeresponsevalid -> dma_subsys_port8:tx_dma_ch1_prefetcher_write_master_writeresponsevalid
	wire  [127:0] dma_subsys_port8_tx_dma_ch1_read_master_readdata;                       // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_read_master_readdata -> dma_subsys_port8:tx_dma_ch1_read_master_readdata
	wire          dma_subsys_port8_tx_dma_ch1_read_master_waitrequest;                    // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_read_master_waitrequest -> dma_subsys_port8:tx_dma_ch1_read_master_waitrequest
	wire   [36:0] dma_subsys_port8_tx_dma_ch1_read_master_address;                        // dma_subsys_port8:tx_dma_ch1_read_master_address -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_read_master_address
	wire          dma_subsys_port8_tx_dma_ch1_read_master_read;                           // dma_subsys_port8:tx_dma_ch1_read_master_read -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_read_master_read
	wire   [15:0] dma_subsys_port8_tx_dma_ch1_read_master_byteenable;                     // dma_subsys_port8:tx_dma_ch1_read_master_byteenable -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_read_master_byteenable
	wire          dma_subsys_port8_tx_dma_ch1_read_master_readdatavalid;                  // mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_read_master_readdatavalid -> dma_subsys_port8:tx_dma_ch1_read_master_readdatavalid
	wire    [4:0] dma_subsys_port8_tx_dma_ch1_read_master_burstcount;                     // dma_subsys_port8:tx_dma_ch1_read_master_burstcount -> mm_interconnect_0:dma_subsys_port8_tx_dma_ch1_read_master_burstcount
	wire  [511:0] mm_interconnect_0_dma_ss_master_s0_readdata;                            // dma_ss_master:s0_readdata -> mm_interconnect_0:dma_ss_master_s0_readdata
	wire          mm_interconnect_0_dma_ss_master_s0_waitrequest;                         // dma_ss_master:s0_waitrequest -> mm_interconnect_0:dma_ss_master_s0_waitrequest
	wire          mm_interconnect_0_dma_ss_master_s0_debugaccess;                         // mm_interconnect_0:dma_ss_master_s0_debugaccess -> dma_ss_master:s0_debugaccess
	wire   [36:0] mm_interconnect_0_dma_ss_master_s0_address;                             // mm_interconnect_0:dma_ss_master_s0_address -> dma_ss_master:s0_address
	wire          mm_interconnect_0_dma_ss_master_s0_read;                                // mm_interconnect_0:dma_ss_master_s0_read -> dma_ss_master:s0_read
	wire   [63:0] mm_interconnect_0_dma_ss_master_s0_byteenable;                          // mm_interconnect_0:dma_ss_master_s0_byteenable -> dma_ss_master:s0_byteenable
	wire          mm_interconnect_0_dma_ss_master_s0_readdatavalid;                       // dma_ss_master:s0_readdatavalid -> mm_interconnect_0:dma_ss_master_s0_readdatavalid
	wire    [1:0] mm_interconnect_0_dma_ss_master_s0_response;                            // dma_ss_master:s0_response -> mm_interconnect_0:dma_ss_master_s0_response
	wire          mm_interconnect_0_dma_ss_master_s0_write;                               // mm_interconnect_0:dma_ss_master_s0_write -> dma_ss_master:s0_write
	wire  [511:0] mm_interconnect_0_dma_ss_master_s0_writedata;                           // mm_interconnect_0:dma_ss_master_s0_writedata -> dma_ss_master:s0_writedata
	wire          mm_interconnect_0_dma_ss_master_s0_writeresponsevalid;                  // dma_ss_master:s0_writeresponsevalid -> mm_interconnect_0:dma_ss_master_s0_writeresponsevalid
	wire    [4:0] mm_interconnect_0_dma_ss_master_s0_burstcount;                          // mm_interconnect_0:dma_ss_master_s0_burstcount -> dma_ss_master:s0_burstcount
	wire          rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> dma_ss_master:reset
	wire          rst_controller_001_reset_out_reset;                                     // rst_controller_001:reset_out -> subsys_ftile_25gbe_1588_dmaclkout_reset:in_reset_n
	wire          rst_controller_002_reset_out_reset;                                     // rst_controller_002:reset_out -> [dma_subsys_port8:rx_dma_resetn, mm_interconnect_0:dma_subsys_port8_rx_dma_resetn_reset_bridge_in_reset_reset]
	wire          rx_dma_reset_bridge_0_out_reset_reset;                                  // rx_dma_reset_bridge_0:out_reset_n -> rst_controller_002:reset_in0
	wire          rst_controller_003_reset_out_reset;                                     // rst_controller_003:reset_out -> dma_subsys_port8:reset_reset_n
	wire          rst_controller_004_reset_out_reset;                                     // rst_controller_004:reset_out -> [mm_interconnect_0:dma_ss_master_reset_reset_bridge_in_reset_reset, mm_interconnect_0:dma_subsys_port8_reset_reset_bridge_in_reset_reset]

	acp_bridge_in_clk acp_bridge_in_clk (
		.in_clk  (iopll_clk_avst_div2_outclk0_clk), //   input,  width = 1,  in_clk.clk
		.out_clk (acp_bridge_in_clk_clk)            //  output,  width = 1, out_clk.clk
	);

	dma_clk_100 dma_clk_100 (
		.in_clk  (dma_clk_100_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (dma_clk_100_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	dma_clk_out_bridge_0 dma_clk_out_bridge_0 (
		.in_clk  (iopll_clk_avst_div2_outclk0_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (dma_clk_out_bridge_0_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	dma_rst_100 dma_rst_100 (
		.clk       (dma_clk_100_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset  (dma_rst_100_in_reset_reset),  //   input,  width = 1,  in_reset.reset
		.out_reset (dma_rst_100_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	dma_ss_master dma_ss_master (
		.clk                   (iopll_clk_avst_div2_outclk0_clk),                       //   input,    width = 1,   clk.clk
		.reset                 (rst_controller_reset_out_reset),                        //   input,    width = 1, reset.reset
		.s0_waitrequest        (mm_interconnect_0_dma_ss_master_s0_waitrequest),        //  output,    width = 1,    s0.waitrequest
		.s0_readdata           (mm_interconnect_0_dma_ss_master_s0_readdata),           //  output,  width = 512,      .readdata
		.s0_readdatavalid      (mm_interconnect_0_dma_ss_master_s0_readdatavalid),      //  output,    width = 1,      .readdatavalid
		.s0_response           (mm_interconnect_0_dma_ss_master_s0_response),           //  output,    width = 2,      .response
		.s0_burstcount         (mm_interconnect_0_dma_ss_master_s0_burstcount),         //   input,    width = 5,      .burstcount
		.s0_writedata          (mm_interconnect_0_dma_ss_master_s0_writedata),          //   input,  width = 512,      .writedata
		.s0_address            (mm_interconnect_0_dma_ss_master_s0_address),            //   input,   width = 37,      .address
		.s0_write              (mm_interconnect_0_dma_ss_master_s0_write),              //   input,    width = 1,      .write
		.s0_read               (mm_interconnect_0_dma_ss_master_s0_read),               //   input,    width = 1,      .read
		.s0_byteenable         (mm_interconnect_0_dma_ss_master_s0_byteenable),         //   input,   width = 64,      .byteenable
		.s0_debugaccess        (mm_interconnect_0_dma_ss_master_s0_debugaccess),        //   input,    width = 1,      .debugaccess
		.s0_writeresponsevalid (mm_interconnect_0_dma_ss_master_s0_writeresponsevalid), //  output,    width = 1,      .writeresponsevalid
		.m0_waitrequest        (dma_ss_master_m0_waitrequest),                          //   input,    width = 1,    m0.waitrequest
		.m0_readdata           (dma_ss_master_m0_readdata),                             //   input,  width = 512,      .readdata
		.m0_readdatavalid      (dma_ss_master_m0_readdatavalid),                        //   input,    width = 1,      .readdatavalid
		.m0_response           (dma_ss_master_m0_response),                             //   input,    width = 2,      .response
		.m0_burstcount         (dma_ss_master_m0_burstcount),                           //  output,    width = 5,      .burstcount
		.m0_writedata          (dma_ss_master_m0_writedata),                            //  output,  width = 512,      .writedata
		.m0_address            (dma_ss_master_m0_address),                              //  output,   width = 37,      .address
		.m0_write              (dma_ss_master_m0_write),                                //  output,    width = 1,      .write
		.m0_read               (dma_ss_master_m0_read),                                 //  output,    width = 1,      .read
		.m0_byteenable         (dma_ss_master_m0_byteenable),                           //  output,   width = 64,      .byteenable
		.m0_debugaccess        (dma_ss_master_m0_debugaccess),                          //  output,    width = 1,      .debugaccess
		.m0_writeresponsevalid (dma_ss_master_m0_writeresponsevalid)                    //   input,    width = 1,      .writeresponsevalid
	);

	ext_hps_m_master ext_hps_m_master (
		.clk                  (dma_clk_100_out_clk_clk),                        //   input,   width = 1,           clock.clk
		.reset                (dma_rst_100_out_reset_reset),                    //   input,   width = 1,           reset.reset
		.avs_s0_address       (ext_hps_m_master_windowed_slave_address),        //   input,  width = 30,  windowed_slave.address
		.avs_s0_read          (ext_hps_m_master_windowed_slave_read),           //   input,   width = 1,                .read
		.avs_s0_readdata      (ext_hps_m_master_windowed_slave_readdata),       //  output,  width = 32,                .readdata
		.avs_s0_write         (ext_hps_m_master_windowed_slave_write),          //   input,   width = 1,                .write
		.avs_s0_writedata     (ext_hps_m_master_windowed_slave_writedata),      //   input,  width = 32,                .writedata
		.avs_s0_readdatavalid (ext_hps_m_master_windowed_slave_readdatavalid),  //  output,   width = 1,                .readdatavalid
		.avs_s0_waitrequest   (ext_hps_m_master_windowed_slave_waitrequest),    //  output,   width = 1,                .waitrequest
		.avs_s0_byteenable    (ext_hps_m_master_windowed_slave_byteenable),     //   input,   width = 4,                .byteenable
		.avs_s0_burstcount    (ext_hps_m_master_windowed_slave_burstcount),     //   input,   width = 1,                .burstcount
		.avm_m0_address       (ext_hps_m_master_expanded_master_address),       //  output,  width = 37, expanded_master.address
		.avm_m0_read          (ext_hps_m_master_expanded_master_read),          //  output,   width = 1,                .read
		.avm_m0_waitrequest   (ext_hps_m_master_expanded_master_waitrequest),   //   input,   width = 1,                .waitrequest
		.avm_m0_readdata      (ext_hps_m_master_expanded_master_readdata),      //   input,  width = 32,                .readdata
		.avm_m0_write         (ext_hps_m_master_expanded_master_write),         //  output,   width = 1,                .write
		.avm_m0_writedata     (ext_hps_m_master_expanded_master_writedata),     //  output,  width = 32,                .writedata
		.avm_m0_readdatavalid (ext_hps_m_master_expanded_master_readdatavalid), //   input,   width = 1,                .readdatavalid
		.avm_m0_byteenable    (ext_hps_m_master_expanded_master_byteenable),    //  output,   width = 4,                .byteenable
		.avm_m0_burstcount    (ext_hps_m_master_expanded_master_burstcount)     //  output,   width = 1,                .burstcount
	);

	iopll_clk_avst_div2 iopll_clk_avst_div2 (
		.rst      (subsys_ftile_25gbe_1588_ninitdone_reset_out_reset_reset), //   input,  width = 1,   reset.reset
		.refclk   (oclk_pll_port8_out_clk_clk),                              //   input,  width = 1,  refclk.clk
		.locked   (),                                                        //  output,  width = 1,  locked.export
		.outclk_0 (iopll_clk_avst_div2_outclk0_clk)                          //  output,  width = 1, outclk0.clk
	);

	oclk_pll_clock_bridge_0 oclk_pll_port8 (
		.in_clk  (oclk_pll_port8_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (oclk_pll_port8_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	rx_dma_reset_bridge_0 rx_dma_reset_bridge_0 (
		.clk         (dma_clk_100_out_clk_clk),                //   input,  width = 1,       clk.clk
		.in_reset_n  (rx_dma_reset_bridge_0_in_reset_reset_n), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (rx_dma_reset_bridge_0_out_reset_reset)   //  output,  width = 1, out_reset.reset_n
	);

	rx_dma_reset_bridge_1 rx_dma_reset_bridge_1 (
		.clk         (dma_clk_100_out_clk_clk),                //   input,  width = 1,       clk.clk
		.in_reset_n  (rx_dma_reset_bridge_1_in_reset_reset_n), //   input,  width = 1,  in_reset.reset_n
		.out_reset_n ()                                        //  output,  width = 1, out_reset.reset_n
	);

	subsys_ftile_25gbe_1588_dmaclkout_reset subsys_ftile_25gbe_1588_dmaclkout_reset (
		.clk         (iopll_clk_avst_div2_outclk0_clk),                           //   input,  width = 1,       clk.clk
		.in_reset_n  (~rst_controller_001_reset_out_reset),                       //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (subsys_ftile_25gbe_1588_dmaclkout_reset_out_reset_reset_n)  //  output,  width = 1, out_reset.reset_n
	);

	subsys_ftile_25gbe_1588_ninitdone_reset subsys_ftile_25gbe_1588_ninitdone_reset (
		.in_reset  (ninit_done_reset),                                        //   input,  width = 1,  in_reset.reset
		.out_reset (subsys_ftile_25gbe_1588_ninitdone_reset_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	subsys_ftile_25gbe_1588 dma_subsys_port8 (
		.rx_dma_resetn                                               (~rst_controller_002_reset_out_reset),                                          //   input,    width = 1,                                   rx_dma_resetn.reset_n
		.csr_waitrequest                                             (dma_subsys_port8_csr_waitrequest),                                             //  output,    width = 1,                                             csr.waitrequest
		.csr_readdata                                                (dma_subsys_port8_csr_readdata),                                                //  output,   width = 32,                                                .readdata
		.csr_readdatavalid                                           (dma_subsys_port8_csr_readdatavalid),                                           //  output,    width = 1,                                                .readdatavalid
		.csr_burstcount                                              (dma_subsys_port8_csr_burstcount),                                              //   input,    width = 1,                                                .burstcount
		.csr_writedata                                               (dma_subsys_port8_csr_writedata),                                               //   input,   width = 32,                                                .writedata
		.csr_address                                                 (dma_subsys_port8_csr_address),                                                 //   input,    width = 8,                                                .address
		.csr_write                                                   (dma_subsys_port8_csr_write),                                                   //   input,    width = 1,                                                .write
		.csr_read                                                    (dma_subsys_port8_csr_read),                                                    //   input,    width = 1,                                                .read
		.csr_byteenable                                              (dma_subsys_port8_csr_byteenable),                                              //   input,    width = 4,                                                .byteenable
		.csr_debugaccess                                             (dma_subsys_port8_csr_debugaccess),                                             //   input,    width = 1,                                                .debugaccess
		.clk_clk                                                     (dma_clk_100_out_clk_clk),                                                      //   input,    width = 1,                                             clk.clk
		.subsys_ftile_25gbe_1588_dmaclkout_in_clk_clk                (iopll_clk_avst_div2_outclk0_clk),                                              //   input,    width = 1,        subsys_ftile_25gbe_1588_dmaclkout_in_clk.clk
		.subsys_ftile_25gbe_1588_o_pll_clk_in_clk_clk                (oclk_pll_port8_out_clk_clk),                                                   //   input,    width = 1,        subsys_ftile_25gbe_1588_o_pll_clk_in_clk.clk
		.reset_reset_n                                               (~rst_controller_003_reset_out_reset),                                          //   input,    width = 1,                                           reset.reset_n
		.ftile_25gbe_rx_dma_ch1_pktin_startofpacket                  (dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_startofpacket),                  //   input,    width = 1,                    ftile_25gbe_rx_dma_ch1_pktin.startofpacket
		.ftile_25gbe_rx_dma_ch1_pktin_valid                          (dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_valid),                          //   input,    width = 1,                                                .valid
		.ftile_25gbe_rx_dma_ch1_pktin_endofpacket                    (dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_endofpacket),                    //   input,    width = 1,                                                .endofpacket
		.ftile_25gbe_rx_dma_ch1_pktin_data                           (dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_data),                           //   input,   width = 64,                                                .data
		.ftile_25gbe_rx_dma_ch1_pktin_empty                          (dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_empty),                          //   input,    width = 3,                                                .empty
		.ftile_25gbe_rx_dma_ch1_pktin_error                          (dma_subsys_port8_ftile_25gbe_rx_dma_ch1_pktin_error),                          //   input,    width = 6,                                                .error
		.ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_valid            (dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_valid),            //   input,    width = 1,      ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts.valid
		.ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_data             (dma_subsys_port8_ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_data),             //   input,   width = 96,                                                .data
		.rx_dma_ch1_prefetcher_read_master_address                   (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_address),                   //  output,   width = 37,               rx_dma_ch1_prefetcher_read_master.address
		.rx_dma_ch1_prefetcher_read_master_read                      (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_read),                      //  output,    width = 1,                                                .read
		.rx_dma_ch1_prefetcher_read_master_readdata                  (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdata),                  //   input,  width = 128,                                                .readdata
		.rx_dma_ch1_prefetcher_read_master_waitrequest               (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_waitrequest),               //   input,    width = 1,                                                .waitrequest
		.rx_dma_ch1_prefetcher_read_master_readdatavalid             (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdatavalid),             //   input,    width = 1,                                                .readdatavalid
		.rx_dma_ch1_prefetcher_read_master_burstcount                (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_burstcount),                //  output,    width = 3,                                                .burstcount
		.rx_dma_ch1_prefetcher_write_master_address                  (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_address),                  //  output,   width = 37,              rx_dma_ch1_prefetcher_write_master.address
		.rx_dma_ch1_prefetcher_write_master_write                    (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_write),                    //  output,    width = 1,                                                .write
		.rx_dma_ch1_prefetcher_write_master_byteenable               (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_byteenable),               //  output,   width = 16,                                                .byteenable
		.rx_dma_ch1_prefetcher_write_master_writedata                (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writedata),                //  output,  width = 128,                                                .writedata
		.rx_dma_ch1_prefetcher_write_master_waitrequest              (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_waitrequest),              //   input,    width = 1,                                                .waitrequest
		.rx_dma_ch1_prefetcher_write_master_response                 (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_response),                 //   input,    width = 2,                                                .response
		.rx_dma_ch1_prefetcher_write_master_writeresponsevalid       (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writeresponsevalid),       //   input,    width = 1,                                                .writeresponsevalid
		.rx_dma_ch1_irq_irq                                          (dma_subsys_port8_rx_dma_ch1_irq_irq),                                          //  output,    width = 1,                                  rx_dma_ch1_irq.irq
		.rx_dma_ch1_write_master_address                             (dma_subsys_port8_rx_dma_ch1_write_master_address),                             //  output,   width = 37,                         rx_dma_ch1_write_master.address
		.rx_dma_ch1_write_master_write                               (dma_subsys_port8_rx_dma_ch1_write_master_write),                               //  output,    width = 1,                                                .write
		.rx_dma_ch1_write_master_byteenable                          (dma_subsys_port8_rx_dma_ch1_write_master_byteenable),                          //  output,   width = 16,                                                .byteenable
		.rx_dma_ch1_write_master_writedata                           (dma_subsys_port8_rx_dma_ch1_write_master_writedata),                           //  output,  width = 128,                                                .writedata
		.rx_dma_ch1_write_master_waitrequest                         (dma_subsys_port8_rx_dma_ch1_write_master_waitrequest),                         //   input,    width = 1,                                                .waitrequest
		.rx_dma_ch1_write_master_burstcount                          (dma_subsys_port8_rx_dma_ch1_write_master_burstcount),                          //  output,    width = 5,                                                .burstcount
		.rx_dma_ch1_write_master_response                            (dma_subsys_port8_rx_dma_ch1_write_master_response),                            //   input,    width = 2,                                                .response
		.rx_dma_ch1_write_master_writeresponsevalid                  (dma_subsys_port8_rx_dma_ch1_write_master_writeresponsevalid),                  //   input,    width = 1,                                                .writeresponsevalid
		.ts_chs_compl_0_clk_bus_in_clk                               (dma_subsys_port8_ts_chs_compl_0_clk_bus_in_clk),                               //   input,    width = 1,                       ts_chs_compl_0_clk_bus_in.clk
		.ts_chs_compl_0_rst_bus_in_reset                             (dma_subsys_port8_ts_chs_compl_0_rst_bus_in_reset),                             //   input,    width = 1,                       ts_chs_compl_0_rst_bus_in.reset
		.ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_valid            (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_valid),            //   input,    width = 1,      ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts.valid
		.ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_fingerprint      (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_fingerprint),      //   input,   width = 20,                                                .fingerprint
		.ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_data             (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_data),             //   input,   width = 96,                                                .data
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready           (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready),           //   input,    width = 1,     ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st.ready
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket   (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket),   //  output,    width = 1,                                                .startofpacket
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid           (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid),           //  output,    width = 1,                                                .valid
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket     (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket),     //  output,    width = 1,                                                .endofpacket
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data            (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data),            //  output,   width = 64,                                                .data
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty           (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty),           //  output,    width = 3,                                                .empty
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error           (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error),           //  output,    width = 1,                                                .error
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_valid       (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_valid),       //  output,    width = 1, ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req.valid
		.ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_fingerprint (dma_subsys_port8_ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_fingerprint), //  output,   width = 20,                                                .fingerprint
		.tx_dma_ch1_prefetcher_read_master_address                   (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_address),                   //  output,   width = 37,               tx_dma_ch1_prefetcher_read_master.address
		.tx_dma_ch1_prefetcher_read_master_read                      (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_read),                      //  output,    width = 1,                                                .read
		.tx_dma_ch1_prefetcher_read_master_readdata                  (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdata),                  //   input,  width = 128,                                                .readdata
		.tx_dma_ch1_prefetcher_read_master_waitrequest               (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_waitrequest),               //   input,    width = 1,                                                .waitrequest
		.tx_dma_ch1_prefetcher_read_master_readdatavalid             (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdatavalid),             //   input,    width = 1,                                                .readdatavalid
		.tx_dma_ch1_prefetcher_read_master_burstcount                (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_burstcount),                //  output,    width = 3,                                                .burstcount
		.tx_dma_ch1_prefetcher_write_master_address                  (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_address),                  //  output,   width = 37,              tx_dma_ch1_prefetcher_write_master.address
		.tx_dma_ch1_prefetcher_write_master_write                    (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_write),                    //  output,    width = 1,                                                .write
		.tx_dma_ch1_prefetcher_write_master_byteenable               (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_byteenable),               //  output,   width = 16,                                                .byteenable
		.tx_dma_ch1_prefetcher_write_master_writedata                (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writedata),                //  output,  width = 128,                                                .writedata
		.tx_dma_ch1_prefetcher_write_master_waitrequest              (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_waitrequest),              //   input,    width = 1,                                                .waitrequest
		.tx_dma_ch1_prefetcher_write_master_response                 (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_response),                 //   input,    width = 2,                                                .response
		.tx_dma_ch1_prefetcher_write_master_writeresponsevalid       (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writeresponsevalid),       //   input,    width = 1,                                                .writeresponsevalid
		.tx_dma_ch1_irq_irq                                          (dma_subsys_port8_tx_dma_ch1_irq_irq),                                          //  output,    width = 1,                                  tx_dma_ch1_irq.irq
		.tx_dma_ch1_read_master_address                              (dma_subsys_port8_tx_dma_ch1_read_master_address),                              //  output,   width = 37,                          tx_dma_ch1_read_master.address
		.tx_dma_ch1_read_master_read                                 (dma_subsys_port8_tx_dma_ch1_read_master_read),                                 //  output,    width = 1,                                                .read
		.tx_dma_ch1_read_master_byteenable                           (dma_subsys_port8_tx_dma_ch1_read_master_byteenable),                           //  output,   width = 16,                                                .byteenable
		.tx_dma_ch1_read_master_readdata                             (dma_subsys_port8_tx_dma_ch1_read_master_readdata),                             //   input,  width = 128,                                                .readdata
		.tx_dma_ch1_read_master_waitrequest                          (dma_subsys_port8_tx_dma_ch1_read_master_waitrequest),                          //   input,    width = 1,                                                .waitrequest
		.tx_dma_ch1_read_master_readdatavalid                        (dma_subsys_port8_tx_dma_ch1_read_master_readdatavalid),                        //   input,    width = 1,                                                .readdatavalid
		.tx_dma_ch1_read_master_burstcount                           (dma_subsys_port8_tx_dma_ch1_read_master_burstcount)                            //  output,    width = 5,                                                .burstcount
	);

	dma_subsystem_altera_mm_interconnect_1920_3nhysga mm_interconnect_0 (
		.dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_address             (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_address),             //   input,   width = 37,   dma_subsys_port8_rx_dma_ch1_prefetcher_read_master.address
		.dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_waitrequest         (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_waitrequest),         //  output,    width = 1,                                                     .waitrequest
		.dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_burstcount          (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_burstcount),          //   input,    width = 3,                                                     .burstcount
		.dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_read                (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_read),                //   input,    width = 1,                                                     .read
		.dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdata            (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdata),            //  output,  width = 128,                                                     .readdata
		.dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdatavalid       (dma_subsys_port8_rx_dma_ch1_prefetcher_read_master_readdatavalid),       //  output,    width = 1,                                                     .readdatavalid
		.dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_address            (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_address),            //   input,   width = 37,  dma_subsys_port8_rx_dma_ch1_prefetcher_write_master.address
		.dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_waitrequest        (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_waitrequest),        //  output,    width = 1,                                                     .waitrequest
		.dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_byteenable         (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_byteenable),         //   input,   width = 16,                                                     .byteenable
		.dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_write              (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_write),              //   input,    width = 1,                                                     .write
		.dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writedata          (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writedata),          //   input,  width = 128,                                                     .writedata
		.dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_response           (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_response),           //  output,    width = 2,                                                     .response
		.dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writeresponsevalid (dma_subsys_port8_rx_dma_ch1_prefetcher_write_master_writeresponsevalid), //  output,    width = 1,                                                     .writeresponsevalid
		.dma_subsys_port8_rx_dma_ch1_write_master_address                       (dma_subsys_port8_rx_dma_ch1_write_master_address),                       //   input,   width = 37,             dma_subsys_port8_rx_dma_ch1_write_master.address
		.dma_subsys_port8_rx_dma_ch1_write_master_waitrequest                   (dma_subsys_port8_rx_dma_ch1_write_master_waitrequest),                   //  output,    width = 1,                                                     .waitrequest
		.dma_subsys_port8_rx_dma_ch1_write_master_burstcount                    (dma_subsys_port8_rx_dma_ch1_write_master_burstcount),                    //   input,    width = 5,                                                     .burstcount
		.dma_subsys_port8_rx_dma_ch1_write_master_byteenable                    (dma_subsys_port8_rx_dma_ch1_write_master_byteenable),                    //   input,   width = 16,                                                     .byteenable
		.dma_subsys_port8_rx_dma_ch1_write_master_write                         (dma_subsys_port8_rx_dma_ch1_write_master_write),                         //   input,    width = 1,                                                     .write
		.dma_subsys_port8_rx_dma_ch1_write_master_writedata                     (dma_subsys_port8_rx_dma_ch1_write_master_writedata),                     //   input,  width = 128,                                                     .writedata
		.dma_subsys_port8_rx_dma_ch1_write_master_response                      (dma_subsys_port8_rx_dma_ch1_write_master_response),                      //  output,    width = 2,                                                     .response
		.dma_subsys_port8_rx_dma_ch1_write_master_writeresponsevalid            (dma_subsys_port8_rx_dma_ch1_write_master_writeresponsevalid),            //  output,    width = 1,                                                     .writeresponsevalid
		.dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_address             (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_address),             //   input,   width = 37,   dma_subsys_port8_tx_dma_ch1_prefetcher_read_master.address
		.dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_waitrequest         (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_waitrequest),         //  output,    width = 1,                                                     .waitrequest
		.dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_burstcount          (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_burstcount),          //   input,    width = 3,                                                     .burstcount
		.dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_read                (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_read),                //   input,    width = 1,                                                     .read
		.dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdata            (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdata),            //  output,  width = 128,                                                     .readdata
		.dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdatavalid       (dma_subsys_port8_tx_dma_ch1_prefetcher_read_master_readdatavalid),       //  output,    width = 1,                                                     .readdatavalid
		.dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_address            (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_address),            //   input,   width = 37,  dma_subsys_port8_tx_dma_ch1_prefetcher_write_master.address
		.dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_waitrequest        (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_waitrequest),        //  output,    width = 1,                                                     .waitrequest
		.dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_byteenable         (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_byteenable),         //   input,   width = 16,                                                     .byteenable
		.dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_write              (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_write),              //   input,    width = 1,                                                     .write
		.dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writedata          (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writedata),          //   input,  width = 128,                                                     .writedata
		.dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_response           (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_response),           //  output,    width = 2,                                                     .response
		.dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writeresponsevalid (dma_subsys_port8_tx_dma_ch1_prefetcher_write_master_writeresponsevalid), //  output,    width = 1,                                                     .writeresponsevalid
		.dma_subsys_port8_tx_dma_ch1_read_master_address                        (dma_subsys_port8_tx_dma_ch1_read_master_address),                        //   input,   width = 37,              dma_subsys_port8_tx_dma_ch1_read_master.address
		.dma_subsys_port8_tx_dma_ch1_read_master_waitrequest                    (dma_subsys_port8_tx_dma_ch1_read_master_waitrequest),                    //  output,    width = 1,                                                     .waitrequest
		.dma_subsys_port8_tx_dma_ch1_read_master_burstcount                     (dma_subsys_port8_tx_dma_ch1_read_master_burstcount),                     //   input,    width = 5,                                                     .burstcount
		.dma_subsys_port8_tx_dma_ch1_read_master_byteenable                     (dma_subsys_port8_tx_dma_ch1_read_master_byteenable),                     //   input,   width = 16,                                                     .byteenable
		.dma_subsys_port8_tx_dma_ch1_read_master_read                           (dma_subsys_port8_tx_dma_ch1_read_master_read),                           //   input,    width = 1,                                                     .read
		.dma_subsys_port8_tx_dma_ch1_read_master_readdata                       (dma_subsys_port8_tx_dma_ch1_read_master_readdata),                       //  output,  width = 128,                                                     .readdata
		.dma_subsys_port8_tx_dma_ch1_read_master_readdatavalid                  (dma_subsys_port8_tx_dma_ch1_read_master_readdatavalid),                  //  output,    width = 1,                                                     .readdatavalid
		.dma_ss_master_s0_address                                               (mm_interconnect_0_dma_ss_master_s0_address),                             //  output,   width = 37,                                     dma_ss_master_s0.address
		.dma_ss_master_s0_write                                                 (mm_interconnect_0_dma_ss_master_s0_write),                               //  output,    width = 1,                                                     .write
		.dma_ss_master_s0_read                                                  (mm_interconnect_0_dma_ss_master_s0_read),                                //  output,    width = 1,                                                     .read
		.dma_ss_master_s0_readdata                                              (mm_interconnect_0_dma_ss_master_s0_readdata),                            //   input,  width = 512,                                                     .readdata
		.dma_ss_master_s0_writedata                                             (mm_interconnect_0_dma_ss_master_s0_writedata),                           //  output,  width = 512,                                                     .writedata
		.dma_ss_master_s0_burstcount                                            (mm_interconnect_0_dma_ss_master_s0_burstcount),                          //  output,    width = 5,                                                     .burstcount
		.dma_ss_master_s0_byteenable                                            (mm_interconnect_0_dma_ss_master_s0_byteenable),                          //  output,   width = 64,                                                     .byteenable
		.dma_ss_master_s0_readdatavalid                                         (mm_interconnect_0_dma_ss_master_s0_readdatavalid),                       //   input,    width = 1,                                                     .readdatavalid
		.dma_ss_master_s0_waitrequest                                           (mm_interconnect_0_dma_ss_master_s0_waitrequest),                         //   input,    width = 1,                                                     .waitrequest
		.dma_ss_master_s0_debugaccess                                           (mm_interconnect_0_dma_ss_master_s0_debugaccess),                         //  output,    width = 1,                                                     .debugaccess
		.dma_ss_master_s0_response                                              (mm_interconnect_0_dma_ss_master_s0_response),                            //   input,    width = 2,                                                     .response
		.dma_ss_master_s0_writeresponsevalid                                    (mm_interconnect_0_dma_ss_master_s0_writeresponsevalid),                  //   input,    width = 1,                                                     .writeresponsevalid
		.dma_subsys_port8_rx_dma_resetn_reset_bridge_in_reset_reset             (rst_controller_002_reset_out_reset),                                     //   input,    width = 1, dma_subsys_port8_rx_dma_resetn_reset_bridge_in_reset.reset
		.dma_subsys_port8_reset_reset_bridge_in_reset_reset                     (rst_controller_004_reset_out_reset),                                     //   input,    width = 1,         dma_subsys_port8_reset_reset_bridge_in_reset.reset
		.dma_ss_master_reset_reset_bridge_in_reset_reset                        (rst_controller_004_reset_out_reset),                                     //   input,    width = 1,            dma_ss_master_reset_reset_bridge_in_reset.reset
		.iopll_clk_avst_div2_outclk0_clk                                        (iopll_clk_avst_div2_outclk0_clk)                                         //   input,    width = 1,                          iopll_clk_avst_div2_outclk0.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (dma_rst_100_out_reset_reset),     //   input,  width = 1, reset_in0.reset
		.clk            (iopll_clk_avst_div2_outclk0_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                // (terminated),                       
		.reset_req_in0  (1'b0),                            // (terminated),                       
		.reset_in1      (1'b0),                            // (terminated),                       
		.reset_req_in1  (1'b0),                            // (terminated),                       
		.reset_in2      (1'b0),                            // (terminated),                       
		.reset_req_in2  (1'b0),                            // (terminated),                       
		.reset_in3      (1'b0),                            // (terminated),                       
		.reset_req_in3  (1'b0),                            // (terminated),                       
		.reset_in4      (1'b0),                            // (terminated),                       
		.reset_req_in4  (1'b0),                            // (terminated),                       
		.reset_in5      (1'b0),                            // (terminated),                       
		.reset_req_in5  (1'b0),                            // (terminated),                       
		.reset_in6      (1'b0),                            // (terminated),                       
		.reset_req_in6  (1'b0),                            // (terminated),                       
		.reset_in7      (1'b0),                            // (terminated),                       
		.reset_req_in7  (1'b0),                            // (terminated),                       
		.reset_in8      (1'b0),                            // (terminated),                       
		.reset_req_in8  (1'b0),                            // (terminated),                       
		.reset_in9      (1'b0),                            // (terminated),                       
		.reset_req_in9  (1'b0),                            // (terminated),                       
		.reset_in10     (1'b0),                            // (terminated),                       
		.reset_req_in10 (1'b0),                            // (terminated),                       
		.reset_in11     (1'b0),                            // (terminated),                       
		.reset_req_in11 (1'b0),                            // (terminated),                       
		.reset_in12     (1'b0),                            // (terminated),                       
		.reset_req_in12 (1'b0),                            // (terminated),                       
		.reset_in13     (1'b0),                            // (terminated),                       
		.reset_req_in13 (1'b0),                            // (terminated),                       
		.reset_in14     (1'b0),                            // (terminated),                       
		.reset_req_in14 (1'b0),                            // (terminated),                       
		.reset_in15     (1'b0),                            // (terminated),                       
		.reset_req_in15 (1'b0)                             // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (subsys_ftile_25gbe_1588_ninitdone_reset_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (iopll_clk_avst_div2_outclk0_clk),                         //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),                      //  output,  width = 1, reset_out.reset
		.reset_req      (),                                                        // (terminated),                       
		.reset_req_in0  (1'b0),                                                    // (terminated),                       
		.reset_in1      (1'b0),                                                    // (terminated),                       
		.reset_req_in1  (1'b0),                                                    // (terminated),                       
		.reset_in2      (1'b0),                                                    // (terminated),                       
		.reset_req_in2  (1'b0),                                                    // (terminated),                       
		.reset_in3      (1'b0),                                                    // (terminated),                       
		.reset_req_in3  (1'b0),                                                    // (terminated),                       
		.reset_in4      (1'b0),                                                    // (terminated),                       
		.reset_req_in4  (1'b0),                                                    // (terminated),                       
		.reset_in5      (1'b0),                                                    // (terminated),                       
		.reset_req_in5  (1'b0),                                                    // (terminated),                       
		.reset_in6      (1'b0),                                                    // (terminated),                       
		.reset_req_in6  (1'b0),                                                    // (terminated),                       
		.reset_in7      (1'b0),                                                    // (terminated),                       
		.reset_req_in7  (1'b0),                                                    // (terminated),                       
		.reset_in8      (1'b0),                                                    // (terminated),                       
		.reset_req_in8  (1'b0),                                                    // (terminated),                       
		.reset_in9      (1'b0),                                                    // (terminated),                       
		.reset_req_in9  (1'b0),                                                    // (terminated),                       
		.reset_in10     (1'b0),                                                    // (terminated),                       
		.reset_req_in10 (1'b0),                                                    // (terminated),                       
		.reset_in11     (1'b0),                                                    // (terminated),                       
		.reset_req_in11 (1'b0),                                                    // (terminated),                       
		.reset_in12     (1'b0),                                                    // (terminated),                       
		.reset_req_in12 (1'b0),                                                    // (terminated),                       
		.reset_in13     (1'b0),                                                    // (terminated),                       
		.reset_req_in13 (1'b0),                                                    // (terminated),                       
		.reset_in14     (1'b0),                                                    // (terminated),                       
		.reset_req_in14 (1'b0),                                                    // (terminated),                       
		.reset_in15     (1'b0),                                                    // (terminated),                       
		.reset_req_in15 (1'b0)                                                     // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~rx_dma_reset_bridge_0_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (iopll_clk_avst_div2_outclk0_clk),        //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (),                                       // (terminated),                       
		.reset_req_in0  (1'b0),                                   // (terminated),                       
		.reset_in1      (1'b0),                                   // (terminated),                       
		.reset_req_in1  (1'b0),                                   // (terminated),                       
		.reset_in2      (1'b0),                                   // (terminated),                       
		.reset_req_in2  (1'b0),                                   // (terminated),                       
		.reset_in3      (1'b0),                                   // (terminated),                       
		.reset_req_in3  (1'b0),                                   // (terminated),                       
		.reset_in4      (1'b0),                                   // (terminated),                       
		.reset_req_in4  (1'b0),                                   // (terminated),                       
		.reset_in5      (1'b0),                                   // (terminated),                       
		.reset_req_in5  (1'b0),                                   // (terminated),                       
		.reset_in6      (1'b0),                                   // (terminated),                       
		.reset_req_in6  (1'b0),                                   // (terminated),                       
		.reset_in7      (1'b0),                                   // (terminated),                       
		.reset_req_in7  (1'b0),                                   // (terminated),                       
		.reset_in8      (1'b0),                                   // (terminated),                       
		.reset_req_in8  (1'b0),                                   // (terminated),                       
		.reset_in9      (1'b0),                                   // (terminated),                       
		.reset_req_in9  (1'b0),                                   // (terminated),                       
		.reset_in10     (1'b0),                                   // (terminated),                       
		.reset_req_in10 (1'b0),                                   // (terminated),                       
		.reset_in11     (1'b0),                                   // (terminated),                       
		.reset_req_in11 (1'b0),                                   // (terminated),                       
		.reset_in12     (1'b0),                                   // (terminated),                       
		.reset_req_in12 (1'b0),                                   // (terminated),                       
		.reset_in13     (1'b0),                                   // (terminated),                       
		.reset_req_in13 (1'b0),                                   // (terminated),                       
		.reset_in14     (1'b0),                                   // (terminated),                       
		.reset_req_in14 (1'b0),                                   // (terminated),                       
		.reset_in15     (1'b0),                                   // (terminated),                       
		.reset_req_in15 (1'b0)                                    // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (dma_rst_100_out_reset_reset),        //   input,  width = 1, reset_in0.reset
		.clk            (dma_clk_100_out_clk_clk),            //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (dma_rst_100_out_reset_reset),        //   input,  width = 1, reset_in0.reset
		.clk            (iopll_clk_avst_div2_outclk0_clk),    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
