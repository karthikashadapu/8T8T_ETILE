// clk_ss.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module clk_ss (
		input  wire  clk_csr_in_clk_clk,                  //                  clk_csr_in_clk.clk
		output wire  clk_csr_out_clk_clk,                 //                 clk_csr_out_clk.clk
		input  wire  clk_dsp_in_clk_clk,                  //                  clk_dsp_in_clk.clk
		output wire  clk_dsp_out_clk_clk,                 //                 clk_dsp_out_clk.clk
		input  wire  clk_eth_in_clk_clk,                  //                  clk_eth_in_clk.clk
		output wire  clk_eth_out_clk_clk,                 //                 clk_eth_out_clk.clk
		input  wire  clk_ftile_402_in_clk_clk,            //            clk_ftile_402_in_clk.clk
		output wire  clk_ftile_402_out_clk_clk,           //           clk_ftile_402_out_clk.clk
		input  wire  clock_bridge_rec_rx_in_clk_clk,      //      clock_bridge_rec_rx_in_clk.clk
		output wire  clock_bridge_rec_rx_out_clk_clk,     //     clock_bridge_rec_rx_out_clk.clk
		output wire  clock_bridge_rec_rx_out_clk_dup_clk, // clock_bridge_rec_rx_out_clk_dup.clk
		input  wire  ftile_in_clk_clk,                    //                    ftile_in_clk.clk
		output wire  ftile_out_clk_clk                    //                   ftile_out_clk.clk
	);

	clk_csr clk_csr (
		.in_clk  (clk_csr_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (clk_csr_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	clk_dsp clk_dsp (
		.in_clk  (clk_dsp_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (clk_dsp_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	clk_eth clk_eth (
		.in_clk  (clk_eth_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (clk_eth_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	clk_ftile_402 clk_ftile_402 (
		.in_clk  (clk_ftile_402_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (clk_ftile_402_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	clk_ss_clock_bridge_rec_rx clk_ss_clock_bridge_rec_rx (
		.in_clk    (clock_bridge_rec_rx_in_clk_clk),      //   input,  width = 1,    in_clk.clk
		.out_clk   (clock_bridge_rec_rx_out_clk_clk),     //  output,  width = 1,   out_clk.clk
		.out_clk_1 (clock_bridge_rec_rx_out_clk_dup_clk)  //  output,  width = 1, out_clk_1.clk
	);

	clk_ss_clock_bridge_0 clock_bridge_0 (
		.in_clk  (ftile_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (ftile_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

endmodule
