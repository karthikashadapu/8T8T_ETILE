// tod_subsys.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module tod_subsys (
		input  wire        cdc_pipeline_0_dst_clk_clk,                              //                             cdc_pipeline_0_dst_clk.clk
		input  wire        cdc_pipeline_0_rst_dst_clk_n_reset_n,                    //                       cdc_pipeline_0_rst_dst_clk_n.reset_n
		output wire [95:0] cdc_pipeline_0_dataout_data,                             //                             cdc_pipeline_0_dataout.data
		input  wire        clock_bridge_100_in_clk_clk,                             //                            clock_bridge_100_in_clk.clk
		input  wire        clock_bridge_156_in_clk_clk,                             //                            clock_bridge_156_in_clk.clk
		input  wire        reset_bridge_100_in_reset_reset_n,                       //                          reset_bridge_100_in_reset.reset_n
		input  wire        reset_bridge_156_in_reset_reset,                         //                          reset_bridge_156_in_reset.reset
		input  wire        tod_timestamp_96b_0_pps_in_pps_in,                       //                         tod_timestamp_96b_0_pps_in.pps_in
		output wire        tod_timestamp_96b_0_rfp_sync_pul_data,                   //                   tod_timestamp_96b_0_rfp_sync_pul.data
		input  wire [4:0]  tod_timestamp_96b_0_tod_timestamp_96b_csr_address,       //          tod_timestamp_96b_0_tod_timestamp_96b_csr.address
		input  wire        tod_timestamp_96b_0_tod_timestamp_96b_csr_write,         //                                                   .write
		input  wire        tod_timestamp_96b_0_tod_timestamp_96b_csr_read,          //                                                   .read
		input  wire [31:0] tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata,     //                                                   .writedata
		output wire [31:0] tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata,      //                                                   .readdata
		output wire        tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest,   //                                                   .waitrequest
		output wire        tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid, //                                                   .readdatavalid
		output wire        tod_timestamp_96b_0_rfp_sync_pul_dup_data,               //               tod_timestamp_96b_0_rfp_sync_pul_dup.data
		input  wire        master_tod_top_0_csr_write,                              //                               master_tod_top_0_csr.write
		input  wire [31:0] master_tod_top_0_csr_writedata,                          //                                                   .writedata
		input  wire        master_tod_top_0_csr_read,                               //                                                   .read
		output wire [31:0] master_tod_top_0_csr_readdata,                           //                                                   .readdata
		output wire        master_tod_top_0_csr_waitrequest,                        //                                                   .waitrequest
		input  wire [3:0]  master_tod_top_0_csr_address,                            //                                                   .address
		input  wire        master_tod_top_0_i_reconfig_rst_n_reset_n,               //                  master_tod_top_0_i_reconfig_rst_n.reset_n
		output wire        master_tod_top_0_pulse_per_second_pps,                   //                  master_tod_top_0_pulse_per_second.pps
		input  wire        mtod_subsys_master_tod_top_0_i_upstr_pll_lock,           //           mtod_subsys_master_tod_top_0_i_upstr_pll.lock
		input  wire        mtod_subsys_clk100_in_clk_clk,                           //                          mtod_subsys_clk100_in_clk.clk
		input  wire        mtod_subsys_pps_load_tod_0_period_clock_clk,             //            mtod_subsys_pps_load_tod_0_period_clock.clk
		input  wire        mtod_subsys_pps_load_tod_0_reset_reset,                  //                   mtod_subsys_pps_load_tod_0_reset.reset
		input  wire        mtod_subsys_pps_load_tod_0_csr_reset_reset,              //               mtod_subsys_pps_load_tod_0_csr_reset.reset
		output wire [31:0] mtod_subsys_pps_load_tod_0_csr_readdata,                 //                     mtod_subsys_pps_load_tod_0_csr.readdata
		input  wire        mtod_subsys_pps_load_tod_0_csr_write,                    //                                                   .write
		input  wire        mtod_subsys_pps_load_tod_0_csr_read,                     //                                                   .read
		input  wire [31:0] mtod_subsys_pps_load_tod_0_csr_writedata,                //                                                   .writedata
		output wire        mtod_subsys_pps_load_tod_0_csr_waitrequest,              //                                                   .waitrequest
		input  wire [5:0]  mtod_subsys_pps_load_tod_0_csr_address,                  //                                                   .address
		input  wire        mtod_subsys_pps_in_pulse_per_second,                     //                                 mtod_subsys_pps_in.pulse_per_second
		output wire        mtod_subsys_pps_load_tod_0_pps_irq_irq,                  //                 mtod_subsys_pps_load_tod_0_pps_irq.irq
		input  wire        mtod_subsys_rstn_in_reset_reset_n,                       //                          mtod_subsys_rstn_in_reset.reset_n
		input  wire        tod_slave_oran_tod_stack_tx_clk_clk,                     //                    tod_slave_oran_tod_stack_tx_clk.clk
		input  wire        tod_slave_oran_tod_stack_rx_clk_clk,                     //                    tod_slave_oran_tod_stack_rx_clk.clk
		input  wire        tod_slave_oran_tod_stack_todsync_sample_clk_clk,         //        tod_slave_oran_tod_stack_todsync_sample_clk.clk
		output wire [95:0] tx_oran_tod_time_of_day_96b_tdata,                       //                        tx_oran_tod_time_of_day_96b.tdata
		output wire        tx_oran_tod_time_of_day_96b_tvalid,                      //                                                   .tvalid
		output wire [95:0] rx_oran_tod_time_of_day_96b_tdata,                       //                        rx_oran_tod_time_of_day_96b.tdata
		output wire        rx_oran_tod_time_of_day_96b_tvalid,                      //                                                   .tvalid
		input  wire        tod_slave_oran_tod_stack_tx_pll_locked_lock,             //             tod_slave_oran_tod_stack_tx_pll_locked.lock
		input  wire        tod_slave_port_8_tod_stack_tx_clk_clk,                   //                  tod_slave_port_8_tod_stack_tx_clk.clk
		input  wire        tod_slave_port_8_tod_stack_rx_clk_clk,                   //                  tod_slave_port_8_tod_stack_rx_clk.clk
		input  wire        tod_slave_port_8_tod_stack_todsync_sample_clk_clk,       //      tod_slave_port_8_tod_stack_todsync_sample_clk.clk
		output wire [95:0] tod_slave_port_8_tod_stack_tx_tod_interface_tdata,       //        tod_slave_port_8_tod_stack_tx_tod_interface.tdata
		output wire        tod_slave_port_8_tod_stack_tx_tod_interface_tvalid,      //                                                   .tvalid
		output wire [95:0] tod_slave_port_8_tod_stack_rx_tod_interface_tdata,       //        tod_slave_port_8_tod_stack_rx_tod_interface.tdata
		output wire        tod_slave_port_8_tod_stack_rx_tod_interface_tvalid,      //                                                   .tvalid
		input  wire        tod_slave_subsys_port_8_tod_stack_tx_pll_locked_lock,    //    tod_slave_subsys_port_8_tod_stack_tx_pll_locked.lock
		input  wire        tod_slave_tod_subsys_clk_100_in_clk_clk,                 //                tod_slave_tod_subsys_clk_100_in_clk.clk
		input  wire        tod_slave_tod_subsys_mtod_clk_in_clk_clk,                //               tod_slave_tod_subsys_mtod_clk_in_clk.clk
		input  wire        tod_slave_tod_subsys_rst_100_in_reset_reset_n,           //              tod_slave_tod_subsys_rst_100_in_reset.reset_n
		input  wire [0:0]  tod_slave_todsync_sample_plllock_split_conduit_end_lock  // tod_slave_todsync_sample_plllock_split_conduit_end.lock
	);

	wire         tod_subsys_clock_bridge_100_out_clk_clk;                     // tod_subsys_clock_bridge_100:out_clk -> [tod_subsys_reset_bridge_100:clk, tod_timestamp_96b_0:clk_100]
	wire         tod_subsys_clock_bridge_156_out_clk_clk;                     // tod_subsys_clock_bridge_156:out_clk -> [cdc_pipeline_0:src_clk, master_tod_subsys_0:master_tod_top_0_i_clk_tod_clk, tod_subsys_reset_bridge_156:clk, tod_sync_interface_adapter_0_0:clk, tod_timestamp_96b_0:clk_tod]
	wire  [95:0] tod_sync_interface_adapter_0_0_tx3_tod_master_data_data;     // tod_sync_interface_adapter_0_0:tx3_tod_master_data -> cdc_pipeline_0:datain
	wire  [95:0] tod_sync_interface_adapter_0_0_tx1_tod_master_data_data;     // tod_sync_interface_adapter_0_0:tx1_tod_master_data -> tod_timestamp_96b_0:eth_tod_master_96b_tx
	wire  [95:0] tod_slave_sub_system_0_master_tod_split_conduit_end_10_data; // tod_slave_sub_system_0:master_tod_split_conduit_end_10_data -> master_tod_subsys_0:mtod_subsys_pps_load_tod_0_time_of_day_96b_data
	wire         master_tod_subsys_0_master_tod_top_0_avst_tod_data_valid;    // master_tod_subsys_0:master_tod_top_0_avst_tod_data_valid -> tod_sync_interface_adapter_0_0:valid
	wire  [95:0] master_tod_subsys_0_master_tod_top_0_avst_tod_data_data;     // master_tod_subsys_0:master_tod_top_0_avst_tod_data_data -> tod_sync_interface_adapter_0_0:time_of_day_96b
	wire         tod_sync_interface_adapter_0_0_tx0_tod_master_data_valid;    // tod_sync_interface_adapter_0_0:valid_0 -> tod_slave_sub_system_0:master_tod_split_conduit_end_valid
	wire  [95:0] tod_sync_interface_adapter_0_0_tx0_tod_master_data_data;     // tod_sync_interface_adapter_0_0:tx0_tod_master_data -> tod_slave_sub_system_0:master_tod_split_conduit_end_data
	wire         tod_subsys_reset_bridge_156_out_reset_reset;                 // tod_subsys_reset_bridge_156:out_reset -> [cdc_pipeline_0:rst_src_clk_n, master_tod_subsys_0:master_tod_top_0_i_tod_rst_n_reset_n, tod_sync_interface_adapter_0_0:rst_n, tod_timestamp_96b_0:rst_clk_tod_n]
	wire         tod_subsys_reset_bridge_100_out_reset_reset;                 // tod_subsys_reset_bridge_100:out_reset_n -> tod_timestamp_96b_0:system_reset_n

	tod_subsys_cdc_pipeline_0 cdc_pipeline_0 (
		.src_clk       (tod_subsys_clock_bridge_156_out_clk_clk),                 //   input,   width = 1,       src_clk.clk
		.rst_src_clk_n (~tod_subsys_reset_bridge_156_out_reset_reset),            //   input,   width = 1, rst_src_clk_n.reset_n
		.dst_clk       (cdc_pipeline_0_dst_clk_clk),                              //   input,   width = 1,       dst_clk.clk
		.rst_dst_clk_n (cdc_pipeline_0_rst_dst_clk_n_reset_n),                    //   input,   width = 1, rst_dst_clk_n.reset_n
		.datain        (tod_sync_interface_adapter_0_0_tx3_tod_master_data_data), //   input,  width = 96,        datain.data
		.dataout       (cdc_pipeline_0_dataout_data)                              //  output,  width = 96,       dataout.data
	);

	tod_subsys_clock_bridge_100 tod_subsys_clock_bridge_100 (
		.in_clk  (clock_bridge_100_in_clk_clk),             //   input,  width = 1,  in_clk.clk
		.out_clk (tod_subsys_clock_bridge_100_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	tod_subsys_clock_bridge_156 tod_subsys_clock_bridge_156 (
		.in_clk  (clock_bridge_156_in_clk_clk),             //   input,  width = 1,  in_clk.clk
		.out_clk (tod_subsys_clock_bridge_156_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	tod_subsys_reset_bridge_100 tod_subsys_reset_bridge_100 (
		.clk         (tod_subsys_clock_bridge_100_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_bridge_100_in_reset_reset_n),           //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (tod_subsys_reset_bridge_100_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	tod_subsys_reset_bridge_156 tod_subsys_reset_bridge_156 (
		.clk       (tod_subsys_clock_bridge_156_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset  (reset_bridge_156_in_reset_reset),             //   input,  width = 1,  in_reset.reset
		.out_reset (tod_subsys_reset_bridge_156_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	tod_subsys_tod_sync_interface_adapter_0_0 tod_sync_interface_adapter_0_0 (
		.time_of_day_96b     (master_tod_subsys_0_master_tod_top_0_avst_tod_data_data),  //   input,  width = 96,     time_of_day_96b.data
		.valid               (master_tod_subsys_0_master_tod_top_0_avst_tod_data_valid), //   input,   width = 1,                    .valid
		.tx0_tod_master_data (tod_sync_interface_adapter_0_0_tx0_tod_master_data_data),  //  output,  width = 96, tx0_tod_master_data.data
		.valid_0             (tod_sync_interface_adapter_0_0_tx0_tod_master_data_valid), //  output,   width = 1,                    .valid
		.tx1_tod_master_data (tod_sync_interface_adapter_0_0_tx1_tod_master_data_data),  //  output,  width = 96, tx1_tod_master_data.data
		.tx2_tod_master_data (),                                                         //  output,  width = 96, tx2_tod_master_data.data
		.tx3_tod_master_data (tod_sync_interface_adapter_0_0_tx3_tod_master_data_data),  //  output,  width = 96, tx3_tod_master_data.data
		.rx0_tod_master_data (),                                                         //  output,  width = 96, rx0_tod_master_data.data
		.clk                 (tod_subsys_clock_bridge_156_out_clk_clk),                  //   input,   width = 1,               clock.clk
		.rst_n               (~tod_subsys_reset_bridge_156_out_reset_reset)              //   input,   width = 1,          reset_sink.reset_n
	);

	tod_subsys_tod_timestamp_96b_0 tod_timestamp_96b_0 (
		.clk_tod                          (tod_subsys_clock_bridge_156_out_clk_clk),                 //   input,    width = 1,                    clk_tod.clk
		.rst_clk_tod_n                    (~tod_subsys_reset_bridge_156_out_reset_reset),            //   input,    width = 1,              rst_clk_tod_n.reset_n
		.clk_100                          (tod_subsys_clock_bridge_100_out_clk_clk),                 //   input,    width = 1,                    clk_100.clk
		.system_reset_n                   (tod_subsys_reset_bridge_100_out_reset_reset),             //   input,    width = 1,             system_reset_n.reset_n
		.pps_in                           (tod_timestamp_96b_0_pps_in_pps_in),                       //   input,    width = 1,                     pps_in.pps_in
		.irq_delay_pulse                  (),                                                        //  output,    width = 1,            irq_delay_pulse.irq
		.eth_tod_master_96b_tx            (tod_sync_interface_adapter_0_0_tx1_tod_master_data_data), //   input,   width = 96,      eth_tod_master_96b_tx.data
		.eth_tod_master_96b_tx_load_data  (),                                                        //  output,   width = 96, eth_tod_master_96b_tx_load.data
		.eth_tod_master_96b_tx_load_valid (),                                                        //  output,    width = 1,                           .valid
		.rfp_sync_pul                     (tod_timestamp_96b_0_rfp_sync_pul_data),                   //  output,    width = 1,               rfp_sync_pul.data
		.rfp_sync_pul_cpri                (),                                                        //  output,    width = 1,          rfp_sync_pul_cpri.cpri_aux_rx_rfp_l1_cpri
		.csr_address                      (tod_timestamp_96b_0_tod_timestamp_96b_csr_address),       //   input,    width = 5,      tod_timestamp_96b_csr.address
		.csr_write                        (tod_timestamp_96b_0_tod_timestamp_96b_csr_write),         //   input,    width = 1,                           .write
		.csr_read                         (tod_timestamp_96b_0_tod_timestamp_96b_csr_read),          //   input,    width = 1,                           .read
		.csr_writedata                    (tod_timestamp_96b_0_tod_timestamp_96b_csr_writedata),     //   input,   width = 32,                           .writedata
		.csr_readdata                     (tod_timestamp_96b_0_tod_timestamp_96b_csr_readdata),      //  output,   width = 32,                           .readdata
		.csr_waitrequest                  (tod_timestamp_96b_0_tod_timestamp_96b_csr_waitrequest),   //  output,    width = 1,                           .waitrequest
		.csr_readdatavalid                (tod_timestamp_96b_0_tod_timestamp_96b_csr_readdatavalid), //  output,    width = 1,                           .readdatavalid
		.ram_read                         (),                                                        //   input,    width = 1,          tod_timestamp_mem.read
		.ram_q                            (),                                                        //  output,  width = 128,                           .readdata
		.rfp_sync_pul_dup                 (tod_timestamp_96b_0_rfp_sync_pul_dup_data)                //  output,    width = 1,           rfp_sync_pul_dup.data
	);

	master_tod_subsys master_tod_subsys_0 (
		.master_tod_top_0_csr_write                                (master_tod_top_0_csr_write),                                  //   input,   width = 1,                       master_tod_top_0_csr.write
		.master_tod_top_0_csr_writedata                            (master_tod_top_0_csr_writedata),                              //   input,  width = 32,                                           .writedata
		.master_tod_top_0_csr_read                                 (master_tod_top_0_csr_read),                                   //   input,   width = 1,                                           .read
		.master_tod_top_0_csr_readdata                             (master_tod_top_0_csr_readdata),                               //  output,  width = 32,                                           .readdata
		.master_tod_top_0_csr_waitrequest                          (master_tod_top_0_csr_waitrequest),                            //  output,   width = 1,                                           .waitrequest
		.master_tod_top_0_csr_address                              (master_tod_top_0_csr_address),                                //   input,   width = 4,                                           .address
		.master_tod_top_0_i_clk_tod_clk                            (tod_subsys_clock_bridge_156_out_clk_clk),                     //   input,   width = 1,                 master_tod_top_0_i_clk_tod.clk
		.master_tod_top_0_i_reconfig_rst_n_reset_n                 (master_tod_top_0_i_reconfig_rst_n_reset_n),                   //   input,   width = 1,          master_tod_top_0_i_reconfig_rst_n.reset_n
		.master_tod_top_0_i_tod_rst_n_reset_n                      (~tod_subsys_reset_bridge_156_out_reset_reset),                //   input,   width = 1,               master_tod_top_0_i_tod_rst_n.reset_n
		.master_tod_top_0_pulse_per_second_pps                     (master_tod_top_0_pulse_per_second_pps),                       //  output,   width = 1,          master_tod_top_0_pulse_per_second.pps
		.master_tod_top_0_avst_tod_data_valid                      (master_tod_subsys_0_master_tod_top_0_avst_tod_data_valid),    //  output,   width = 1,             master_tod_top_0_avst_tod_data.valid
		.master_tod_top_0_avst_tod_data_data                       (master_tod_subsys_0_master_tod_top_0_avst_tod_data_data),     //  output,  width = 96,                                           .data
		.master_tod_top_0_i_upstr_pll_lock                         (mtod_subsys_master_tod_top_0_i_upstr_pll_lock),               //   input,   width = 1,               master_tod_top_0_i_upstr_pll.lock
		.mtod_subsys_clk100_in_clk_clk                             (mtod_subsys_clk100_in_clk_clk),                               //   input,   width = 1,                  mtod_subsys_clk100_in_clk.clk
		.mtod_subsys_pps_load_tod_0_period_clock_clk               (mtod_subsys_pps_load_tod_0_period_clock_clk),                 //   input,   width = 1,    mtod_subsys_pps_load_tod_0_period_clock.clk
		.mtod_subsys_pps_load_tod_0_reset_reset                    (mtod_subsys_pps_load_tod_0_reset_reset),                      //   input,   width = 1,           mtod_subsys_pps_load_tod_0_reset.reset
		.mtod_subsys_pps_load_tod_0_csr_reset_reset                (mtod_subsys_pps_load_tod_0_csr_reset_reset),                  //   input,   width = 1,       mtod_subsys_pps_load_tod_0_csr_reset.reset
		.mtod_subsys_pps_load_tod_0_csr_readdata                   (mtod_subsys_pps_load_tod_0_csr_readdata),                     //  output,  width = 32,             mtod_subsys_pps_load_tod_0_csr.readdata
		.mtod_subsys_pps_load_tod_0_csr_write                      (mtod_subsys_pps_load_tod_0_csr_write),                        //   input,   width = 1,                                           .write
		.mtod_subsys_pps_load_tod_0_csr_read                       (mtod_subsys_pps_load_tod_0_csr_read),                         //   input,   width = 1,                                           .read
		.mtod_subsys_pps_load_tod_0_csr_writedata                  (mtod_subsys_pps_load_tod_0_csr_writedata),                    //   input,  width = 32,                                           .writedata
		.mtod_subsys_pps_load_tod_0_csr_waitrequest                (mtod_subsys_pps_load_tod_0_csr_waitrequest),                  //  output,   width = 1,                                           .waitrequest
		.mtod_subsys_pps_load_tod_0_csr_address                    (mtod_subsys_pps_load_tod_0_csr_address),                      //   input,   width = 6,                                           .address
		.mtod_subsys_pps_load_tod_0_pps_interface_pulse_per_second (mtod_subsys_pps_in_pulse_per_second),                         //   input,   width = 1,   mtod_subsys_pps_load_tod_0_pps_interface.pulse_per_second
		.mtod_subsys_pps_load_tod_0_time_of_day_96b_data           (tod_slave_sub_system_0_master_tod_split_conduit_end_10_data), //   input,  width = 96, mtod_subsys_pps_load_tod_0_time_of_day_96b.data
		.mtod_subsys_pps_load_tod_0_pps_irq_irq                    (mtod_subsys_pps_load_tod_0_pps_irq_irq),                      //  output,   width = 1,         mtod_subsys_pps_load_tod_0_pps_irq.irq
		.mtod_subsys_rstn_in_reset_reset_n                         (mtod_subsys_rstn_in_reset_reset_n)                            //   input,   width = 1,                  mtod_subsys_rstn_in_reset.reset_n
	);

	tod_slave_sub_system tod_slave_sub_system_0 (
		.master_tod_split_conduit_end_data             (tod_sync_interface_adapter_0_0_tx0_tod_master_data_data),     //   input,  width = 96,             master_tod_split_conduit_end.data
		.master_tod_split_conduit_end_valid            (tod_sync_interface_adapter_0_0_tx0_tod_master_data_valid),    //   input,   width = 1,                                         .valid
		.master_tod_split_conduit_end_10_data          (tod_slave_sub_system_0_master_tod_split_conduit_end_10_data), //  output,  width = 96,          master_tod_split_conduit_end_10.data
		.master_tod_split_conduit_end_10_valid         (),                                                            //  output,   width = 1,                                         .valid
		.oran_tod_stack_tx_clk_clk                     (tod_slave_oran_tod_stack_tx_clk_clk),                         //   input,   width = 1,                    oran_tod_stack_tx_clk.clk
		.oran_tod_stack_rx_clk_clk                     (tod_slave_oran_tod_stack_rx_clk_clk),                         //   input,   width = 1,                    oran_tod_stack_rx_clk.clk
		.oran_tod_stack_todsync_sample_clk_clk         (tod_slave_oran_tod_stack_todsync_sample_clk_clk),             //   input,   width = 1,        oran_tod_stack_todsync_sample_clk.clk
		.oran_tod_stack_tx_tod_interface_tdata         (tx_oran_tod_time_of_day_96b_tdata),                           //  output,  width = 96,          oran_tod_stack_tx_tod_interface.tdata
		.oran_tod_stack_tx_tod_interface_tvalid        (tx_oran_tod_time_of_day_96b_tvalid),                          //  output,   width = 1,                                         .tvalid
		.oran_tod_stack_rx_tod_interface_tdata         (rx_oran_tod_time_of_day_96b_tdata),                           //  output,  width = 96,          oran_tod_stack_rx_tod_interface.tdata
		.oran_tod_stack_rx_tod_interface_tvalid        (rx_oran_tod_time_of_day_96b_tvalid),                          //  output,   width = 1,                                         .tvalid
		.oran_tod_stack_tx_pll_locked_lock             (tod_slave_oran_tod_stack_tx_pll_locked_lock),                 //   input,   width = 1,             oran_tod_stack_tx_pll_locked.lock
		.port_8_tod_stack_tx_clk_clk                   (tod_slave_port_8_tod_stack_tx_clk_clk),                       //   input,   width = 1,                  port_8_tod_stack_tx_clk.clk
		.port_8_tod_stack_rx_clk_clk                   (tod_slave_port_8_tod_stack_rx_clk_clk),                       //   input,   width = 1,                  port_8_tod_stack_rx_clk.clk
		.port_8_tod_stack_todsync_sample_clk_clk       (tod_slave_port_8_tod_stack_todsync_sample_clk_clk),           //   input,   width = 1,      port_8_tod_stack_todsync_sample_clk.clk
		.port_8_tod_stack_tx_tod_interface_tdata       (tod_slave_port_8_tod_stack_tx_tod_interface_tdata),           //  output,  width = 96,        port_8_tod_stack_tx_tod_interface.tdata
		.port_8_tod_stack_tx_tod_interface_tvalid      (tod_slave_port_8_tod_stack_tx_tod_interface_tvalid),          //  output,   width = 1,                                         .tvalid
		.port_8_tod_stack_rx_tod_interface_tdata       (tod_slave_port_8_tod_stack_rx_tod_interface_tdata),           //  output,  width = 96,        port_8_tod_stack_rx_tod_interface.tdata
		.port_8_tod_stack_rx_tod_interface_tvalid      (tod_slave_port_8_tod_stack_rx_tod_interface_tvalid),          //  output,   width = 1,                                         .tvalid
		.port_8_tod_stack_tx_pll_locked_lock           (tod_slave_subsys_port_8_tod_stack_tx_pll_locked_lock),        //   input,   width = 1,           port_8_tod_stack_tx_pll_locked.lock
		.tod_subsys_clk_100_in_clk_clk                 (tod_slave_tod_subsys_clk_100_in_clk_clk),                     //   input,   width = 1,                tod_subsys_clk_100_in_clk.clk
		.tod_subsys_mtod_clk_in_clk_clk                (tod_slave_tod_subsys_mtod_clk_in_clk_clk),                    //   input,   width = 1,               tod_subsys_mtod_clk_in_clk.clk
		.tod_subsys_rst_100_in_reset_reset_n           (tod_slave_tod_subsys_rst_100_in_reset_reset_n),               //   input,   width = 1,              tod_subsys_rst_100_in_reset.reset_n
		.todsync_sample_plllock_split_conduit_end_lock (tod_slave_todsync_sample_plllock_split_conduit_end_lock)      //   input,   width = 1, todsync_sample_plllock_split_conduit_end.lock
	);

endmodule
