// oran_tod_subsys.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module oran_tod_subsys (
		input  wire        eth_1588_tod_synchronizer_clk_master_clk,      //     eth_1588_tod_synchronizer_clk_master.clk
		input  wire        eth_1588_tod_synchronizer_reset_master_reset,  //   eth_1588_tod_synchronizer_reset_master.reset
		input  wire        eth_1588_tod_synchronizer_clk_slave_clk,       //      eth_1588_tod_synchronizer_clk_slave.clk
		input  wire        eth_1588_tod_synchronizer_reset_slave_reset,   //    eth_1588_tod_synchronizer_reset_slave.reset
		input  wire        eth_1588_tod_synchronizer_clk_sampling_clk,    //   eth_1588_tod_synchronizer_clk_sampling.clk
		input  wire        eth_1588_tod_synchronizer_start_tod_sync_data, // eth_1588_tod_synchronizer_start_tod_sync.data
		output wire [95:0] oran_tod_time_of_day_96b_data,                 //                 oran_tod_time_of_day_96b.data
		output wire        oran_tod_time_of_day_96b_valid,                //                                         .valid
		input  wire        rst_tod_n_reset_n,                             //                                rst_tod_n.reset_n
		input  wire [95:0] ptp_seconds_data,                              //                              ptp_seconds.data
		input  wire        clk_tod_clk                                    //                                  clk_tod.clk
	);

	wire  [95:0] ptp2gps_conv_0_gps_seconds_data; // ptp2gps_conv_0:gps_seconds -> eth_1588_tod_synchronizer:tod_master_data

	eth_1588_tod_synchronizer eth_1588_tod_synchronizer (
		.clk_master      (eth_1588_tod_synchronizer_clk_master_clk),      //   input,   width = 1,      clk_master.clk
		.reset_master    (eth_1588_tod_synchronizer_reset_master_reset),  //   input,   width = 1,    reset_master.reset
		.clk_slave       (eth_1588_tod_synchronizer_clk_slave_clk),       //   input,   width = 1,       clk_slave.clk
		.reset_slave     (eth_1588_tod_synchronizer_reset_slave_reset),   //   input,   width = 1,     reset_slave.reset
		.clk_sampling    (eth_1588_tod_synchronizer_clk_sampling_clk),    //   input,   width = 1,    clk_sampling.clk
		.start_tod_sync  (eth_1588_tod_synchronizer_start_tod_sync_data), //   input,   width = 1,  start_tod_sync.data
		.tod_master_data (ptp2gps_conv_0_gps_seconds_data),               //   input,  width = 96, tod_master_data.data
		.tod_slave_data  (oran_tod_time_of_day_96b_data),                 //  output,  width = 96,  tod_slave_data.data
		.tod_slave_valid (oran_tod_time_of_day_96b_valid)                 //  output,   width = 1,                .valid
	);

	oran_tod_subsys_ptp2gps_conv_0 ptp2gps_conv_0 (
		.rst_tod_n   (rst_tod_n_reset_n),               //   input,   width = 1,   rst_tod_n.reset_n
		.ptp_seconds (ptp_seconds_data),                //   input,  width = 96, ptp_seconds.data
		.gps_seconds (ptp2gps_conv_0_gps_seconds_data), //  output,  width = 96, gps_seconds.data
		.clk_tod     (clk_tod_clk)                      //   input,   width = 1,     clk_tod.clk
	);

endmodule
