// ed_synth.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module ed_synth (
		input  wire         capture_if_reset_soft_n_rst_soft_n,                 //        capture_if_reset_soft_n.rst_soft_n
		input  wire [55:0]  capture_if_radio_config_status_radio_config_status, // capture_if_radio_config_status.radio_config_status
		input  wire         lphy_avst_sink_dsp_capture_valid,                   //     lphy_avst_sink_dsp_capture.valid
		input  wire [31:0]  lphy_avst_sink_dsp_capture_data,                    //                               .data
		input  wire [2:0]   lphy_avst_sink_dsp_capture_channel,                 //                               .channel
		input  wire         dxc_avst_sink_dsp_capture_valid,                    //      dxc_avst_sink_dsp_capture.valid
		input  wire [31:0]  dxc_avst_sink_dsp_capture_data,                     //                               .data
		input  wire [2:0]   dxc_avst_sink_dsp_capture_channel,                  //                               .channel
		output wire [31:0]  interface_sel_data,                                 //                  interface_sel.data
		input  wire         dsp_in_clk_clk,                                     //                     dsp_in_clk.clk
		input  wire         eth_in_clk_clk,                                     //                     eth_in_clk.clk
		input  wire         clock_csr_clk,                                      //                      clock_csr.clk
		input  wire         clock_bridge_dspby2_in_clk_clk,                     //     clock_bridge_dspby2_in_clk.clk
		output wire         ed_synth_h2f_bridge_s0_waitrequest,                 //         ed_synth_h2f_bridge_s0.waitrequest
		output wire [511:0] ed_synth_h2f_bridge_s0_readdata,                    //                               .readdata
		output wire         ed_synth_h2f_bridge_s0_readdatavalid,               //                               .readdatavalid
		input  wire [0:0]   ed_synth_h2f_bridge_s0_burstcount,                  //                               .burstcount
		input  wire [511:0] ed_synth_h2f_bridge_s0_writedata,                   //                               .writedata
		input  wire [27:0]  ed_synth_h2f_bridge_s0_address,                     //                               .address
		input  wire         ed_synth_h2f_bridge_s0_write,                       //                               .write
		input  wire         ed_synth_h2f_bridge_s0_read,                        //                               .read
		input  wire [63:0]  ed_synth_h2f_bridge_s0_byteenable,                  //                               .byteenable
		input  wire         ed_synth_h2f_bridge_s0_debugaccess,                 //                               .debugaccess
		output wire         h2f_lw_bridge_s0_waitrequest,                       //               h2f_lw_bridge_s0.waitrequest
		output wire [31:0]  h2f_lw_bridge_s0_readdata,                          //                               .readdata
		output wire         h2f_lw_bridge_s0_readdatavalid,                     //                               .readdatavalid
		input  wire [0:0]   h2f_lw_bridge_s0_burstcount,                        //                               .burstcount
		input  wire [31:0]  h2f_lw_bridge_s0_writedata,                         //                               .writedata
		input  wire [12:0]  h2f_lw_bridge_s0_address,                           //                               .address
		input  wire         h2f_lw_bridge_s0_write,                             //                               .write
		input  wire         h2f_lw_bridge_s0_read,                              //                               .read
		input  wire [3:0]   h2f_lw_bridge_s0_byteenable,                        //                               .byteenable
		input  wire         h2f_lw_bridge_s0_debugaccess,                       //                               .debugaccess
		input  wire         dsp_in_reset_reset_n,                               //                   dsp_in_reset.reset_n
		input  wire         eth_in_reset_reset_n,                               //                   eth_in_reset.reset_n
		input  wire         reset_csr_reset_n,                                  //                      reset_csr.reset_n
		output wire         wr_msgdma_0_csr_irq_irq                             //            wr_msgdma_0_csr_irq.irq
	);

	wire          capture_if_top_0_avst_source_capture_valid;                       // capture_if_top_0:avst_src_capture_valid -> ddr4_wr_rd_0:wr_msgdma_0_st_sink_valid
	wire  [127:0] capture_if_top_0_avst_source_capture_data;                        // capture_if_top_0:avst_src_capture_data -> ddr4_wr_rd_0:wr_msgdma_0_st_sink_data
	wire          capture_if_top_0_avst_source_capture_ready;                       // ddr4_wr_rd_0:wr_msgdma_0_st_sink_ready -> capture_if_top_0:avst_src_capture_ready
	wire          clock_csr_out_clk_clk;                                            // clock_csr:out_clk -> [capture_if_top_0:clk_csr, ddr4_wr_rd_0:ocm_rd_clk_clk, ed_synth_h2f_bridge:clk, ed_synth_h2f_lw_bridge:clk, mm_interconnect_0:clock_csr_out_clk_clk, mm_interconnect_1:clock_csr_out_clk_clk, reset_csr:clk, rst_controller:clk, rst_controller_002:clk]
	wire          clock_bridge_dsp_out_clk_clk;                                     // clock_bridge_dsp:out_clk -> [capture_if_top_0:clk_dsp, ed_synth_reset_bridge_dsp:clk]
	wire          clock_bridge_eth_out_clk_clk;                                     // clock_bridge_eth:out_clk -> [capture_if_top_0:clk_eth_xran_ul, ed_synth_reset_bridge_eth:clk]
	wire          ed_synth_clock_bridge_dspby2_out_clk_clk;                         // ed_synth_clock_bridge_dspby2:out_clk -> [capture_if_top_0:clk_capture_dma, ddr4_wr_rd_0:in_clk_clk, mm_interconnect_0:ed_synth_clock_bridge_dspby2_out_clk_clk, mm_interconnect_1:ed_synth_clock_bridge_dspby2_out_clk_clk, rst_controller_001:clk, rst_controller_003:clk]
	wire          ed_synth_reset_bridge_dsp_out_reset_reset;                        // ed_synth_reset_bridge_dsp:out_reset_n -> capture_if_top_0:rst_dsp_n
	wire          ed_synth_reset_bridge_eth_out_reset_reset;                        // ed_synth_reset_bridge_eth:out_reset_n -> capture_if_top_0:rst_eth_xran_n_ul
	wire          ed_synth_h2f_lw_bridge_m0_waitrequest;                            // mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_waitrequest -> ed_synth_h2f_lw_bridge:m0_waitrequest
	wire   [31:0] ed_synth_h2f_lw_bridge_m0_readdata;                               // mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_readdata -> ed_synth_h2f_lw_bridge:m0_readdata
	wire          ed_synth_h2f_lw_bridge_m0_debugaccess;                            // ed_synth_h2f_lw_bridge:m0_debugaccess -> mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_debugaccess
	wire   [12:0] ed_synth_h2f_lw_bridge_m0_address;                                // ed_synth_h2f_lw_bridge:m0_address -> mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_address
	wire          ed_synth_h2f_lw_bridge_m0_read;                                   // ed_synth_h2f_lw_bridge:m0_read -> mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_read
	wire    [3:0] ed_synth_h2f_lw_bridge_m0_byteenable;                             // ed_synth_h2f_lw_bridge:m0_byteenable -> mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_byteenable
	wire          ed_synth_h2f_lw_bridge_m0_readdatavalid;                          // mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_readdatavalid -> ed_synth_h2f_lw_bridge:m0_readdatavalid
	wire   [31:0] ed_synth_h2f_lw_bridge_m0_writedata;                              // ed_synth_h2f_lw_bridge:m0_writedata -> mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_writedata
	wire          ed_synth_h2f_lw_bridge_m0_write;                                  // ed_synth_h2f_lw_bridge:m0_write -> mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_write
	wire    [0:0] ed_synth_h2f_lw_bridge_m0_burstcount;                             // ed_synth_h2f_lw_bridge:m0_burstcount -> mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_burstcount
	wire   [31:0] mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_readdata;            // ddr4_wr_rd_0:csr_bridge_s0_readdata -> mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_readdata
	wire          mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_waitrequest;         // ddr4_wr_rd_0:csr_bridge_s0_waitrequest -> mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_waitrequest
	wire          mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_debugaccess;         // mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_debugaccess -> ddr4_wr_rd_0:csr_bridge_s0_debugaccess
	wire    [5:0] mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_address;             // mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_address -> ddr4_wr_rd_0:csr_bridge_s0_address
	wire          mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_read;                // mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_read -> ddr4_wr_rd_0:csr_bridge_s0_read
	wire    [3:0] mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_byteenable;          // mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_byteenable -> ddr4_wr_rd_0:csr_bridge_s0_byteenable
	wire          mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_readdatavalid;       // ddr4_wr_rd_0:csr_bridge_s0_readdatavalid -> mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_readdatavalid
	wire          mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_write;               // mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_write -> ddr4_wr_rd_0:csr_bridge_s0_write
	wire   [31:0] mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_writedata;           // mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_writedata -> ddr4_wr_rd_0:csr_bridge_s0_writedata
	wire    [0:0] mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_burstcount;          // mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_burstcount -> ddr4_wr_rd_0:csr_bridge_s0_burstcount
	wire   [31:0] mm_interconnect_0_capture_if_top_0_csr_dsp_capture_readdata;      // capture_if_top_0:csr_dsp_capture_readdata -> mm_interconnect_0:capture_if_top_0_csr_dsp_capture_readdata
	wire          mm_interconnect_0_capture_if_top_0_csr_dsp_capture_waitrequest;   // capture_if_top_0:csr_dsp_capture_waitrequest -> mm_interconnect_0:capture_if_top_0_csr_dsp_capture_waitrequest
	wire    [4:0] mm_interconnect_0_capture_if_top_0_csr_dsp_capture_address;       // mm_interconnect_0:capture_if_top_0_csr_dsp_capture_address -> capture_if_top_0:csr_dsp_capture_address
	wire          mm_interconnect_0_capture_if_top_0_csr_dsp_capture_read;          // mm_interconnect_0:capture_if_top_0_csr_dsp_capture_read -> capture_if_top_0:csr_dsp_capture_read
	wire          mm_interconnect_0_capture_if_top_0_csr_dsp_capture_readdatavalid; // capture_if_top_0:csr_dsp_capture_readdatavalid -> mm_interconnect_0:capture_if_top_0_csr_dsp_capture_readdatavalid
	wire          mm_interconnect_0_capture_if_top_0_csr_dsp_capture_write;         // mm_interconnect_0:capture_if_top_0_csr_dsp_capture_write -> capture_if_top_0:csr_dsp_capture_write
	wire   [31:0] mm_interconnect_0_capture_if_top_0_csr_dsp_capture_writedata;     // mm_interconnect_0:capture_if_top_0_csr_dsp_capture_writedata -> capture_if_top_0:csr_dsp_capture_writedata
	wire          ed_synth_h2f_bridge_m0_waitrequest;                               // mm_interconnect_1:ed_synth_h2f_bridge_m0_waitrequest -> ed_synth_h2f_bridge:m0_waitrequest
	wire  [511:0] ed_synth_h2f_bridge_m0_readdata;                                  // mm_interconnect_1:ed_synth_h2f_bridge_m0_readdata -> ed_synth_h2f_bridge:m0_readdata
	wire          ed_synth_h2f_bridge_m0_debugaccess;                               // ed_synth_h2f_bridge:m0_debugaccess -> mm_interconnect_1:ed_synth_h2f_bridge_m0_debugaccess
	wire   [27:0] ed_synth_h2f_bridge_m0_address;                                   // ed_synth_h2f_bridge:m0_address -> mm_interconnect_1:ed_synth_h2f_bridge_m0_address
	wire          ed_synth_h2f_bridge_m0_read;                                      // ed_synth_h2f_bridge:m0_read -> mm_interconnect_1:ed_synth_h2f_bridge_m0_read
	wire   [63:0] ed_synth_h2f_bridge_m0_byteenable;                                // ed_synth_h2f_bridge:m0_byteenable -> mm_interconnect_1:ed_synth_h2f_bridge_m0_byteenable
	wire          ed_synth_h2f_bridge_m0_readdatavalid;                             // mm_interconnect_1:ed_synth_h2f_bridge_m0_readdatavalid -> ed_synth_h2f_bridge:m0_readdatavalid
	wire  [511:0] ed_synth_h2f_bridge_m0_writedata;                                 // ed_synth_h2f_bridge:m0_writedata -> mm_interconnect_1:ed_synth_h2f_bridge_m0_writedata
	wire          ed_synth_h2f_bridge_m0_write;                                     // ed_synth_h2f_bridge:m0_write -> mm_interconnect_1:ed_synth_h2f_bridge_m0_write
	wire    [0:0] ed_synth_h2f_bridge_m0_burstcount;                                // ed_synth_h2f_bridge:m0_burstcount -> mm_interconnect_1:ed_synth_h2f_bridge_m0_burstcount
	wire  [127:0] mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_readdata;          // ddr4_wr_rd_0:emif_mm_slave_1_readdata -> mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_readdata
	wire          mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_waitrequest;       // ddr4_wr_rd_0:emif_mm_slave_1_waitrequest -> mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_waitrequest
	wire   [20:0] mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_address;           // mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_address -> ddr4_wr_rd_0:emif_mm_slave_1_address
	wire          mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_read;              // mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_read -> ddr4_wr_rd_0:emif_mm_slave_1_read
	wire   [15:0] mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_byteenable;        // mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_byteenable -> ddr4_wr_rd_0:emif_mm_slave_1_byteenable
	wire          mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_readdatavalid;     // ddr4_wr_rd_0:emif_mm_slave_1_readdatavalid -> mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_readdatavalid
	wire          mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_write;             // mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_write -> ddr4_wr_rd_0:emif_mm_slave_1_write
	wire  [127:0] mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_writedata;         // mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_writedata -> ddr4_wr_rd_0:emif_mm_slave_1_writedata
	wire    [6:0] mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_burstcount;        // mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_burstcount -> ddr4_wr_rd_0:emif_mm_slave_1_burstcount
	wire  [127:0] mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_readdata;                   // ddr4_wr_rd_0:ocm_rd_readdata -> mm_interconnect_1:ddr4_wr_rd_0_ocm_rd_readdata
	wire   [12:0] mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_address;                    // mm_interconnect_1:ddr4_wr_rd_0_ocm_rd_address -> ddr4_wr_rd_0:ocm_rd_address
	wire          mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_read;                       // mm_interconnect_1:ddr4_wr_rd_0_ocm_rd_read -> ddr4_wr_rd_0:ocm_rd_read
	wire          rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [capture_if_top_0:rst_csr_n, ddr4_wr_rd_0:ocm_rd_reset_reset, ed_synth_h2f_bridge:reset, ed_synth_h2f_lw_bridge:reset, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [ddr4_wr_rd_0:ocm_rd_reset_reset_req, rst_translator:reset_req_in]
	wire          reset_csr_out_reset_reset;                                        // reset_csr:out_reset_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	wire          rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [capture_if_top_0:rst_capture_dma_n, ddr4_wr_rd_0:in_reset_reset_n]
	wire          rst_controller_002_reset_out_reset;                               // rst_controller_002:reset_out -> [mm_interconnect_0:ed_synth_h2f_lw_bridge_m0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:ed_synth_h2f_lw_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ed_synth_h2f_bridge_m0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ed_synth_h2f_bridge_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                               // rst_controller_003:reset_out -> [mm_interconnect_0:ddr4_wr_rd_0_csr_bridge_s0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:ddr4_wr_rd_0_in_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ddr4_wr_rd_0_emif_mm_slave_1_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ddr4_wr_rd_0_in_reset_reset_bridge_in_reset_reset]

	ed_synth_capture_if_top_0 capture_if_top_0 (
		.csr_dsp_capture_address          (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_address),       //   input,    width = 5,            csr_dsp_capture.address
		.csr_dsp_capture_write            (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_write),         //   input,    width = 1,                           .write
		.csr_dsp_capture_read             (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_read),          //   input,    width = 1,                           .read
		.csr_dsp_capture_writedata        (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_writedata),     //   input,   width = 32,                           .writedata
		.csr_dsp_capture_readdata         (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_readdata),      //  output,   width = 32,                           .readdata
		.csr_dsp_capture_waitrequest      (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_waitrequest),   //  output,    width = 1,                           .waitrequest
		.csr_dsp_capture_readdatavalid    (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_readdatavalid), //  output,    width = 1,                           .readdatavalid
		.clk_dsp                          (clock_bridge_dsp_out_clk_clk),                                     //   input,    width = 1,                  clock_dsp.clk
		.clk_csr                          (clock_csr_out_clk_clk),                                            //   input,    width = 1,                  clock_csr.clk
		.clk_eth_xran_ul                  (clock_bridge_eth_out_clk_clk),                                     //   input,    width = 1,                  clock_eth.clk
		.clk_capture_dma                  (ed_synth_clock_bridge_dspby2_out_clk_clk),                         //   input,    width = 1,                  clock_dma.clk
		.rst_csr_n                        (~rst_controller_reset_out_reset),                                  //   input,    width = 1,                reset_csr_n.reset_n
		.rst_dsp_n                        (ed_synth_reset_bridge_dsp_out_reset_reset),                        //   input,    width = 1,                reset_dsp_n.reset_n
		.rst_eth_xran_n_ul                (ed_synth_reset_bridge_eth_out_reset_reset),                        //   input,    width = 1,                reset_eth_n.reset_n
		.rst_capture_dma_n                (~rst_controller_001_reset_out_reset),                              //   input,    width = 1,                reset_dma_n.reset_n
		.rst_soft_n                       (capture_if_reset_soft_n_rst_soft_n),                               //   input,    width = 1,               reset_soft_n.rst_soft_n
		.avst_src_capture_valid           (capture_if_top_0_avst_source_capture_valid),                       //  output,    width = 1,        avst_source_capture.valid
		.avst_src_capture_data            (capture_if_top_0_avst_source_capture_data),                        //  output,  width = 128,                           .data
		.avst_src_capture_ready           (capture_if_top_0_avst_source_capture_ready),                       //   input,    width = 1,                           .ready
		.radio_config_status              (capture_if_radio_config_status_radio_config_status),               //   input,   width = 56,        radio_config_status.radio_config_status
		.lphy_avst_sink_dsp_capture_valid (lphy_avst_sink_dsp_capture_valid),                                 //   input,    width = 1, lphy_avst_sink_dsp_capture.valid
		.lphy_avst_sink_dsp_capture_data  (lphy_avst_sink_dsp_capture_data),                                  //   input,   width = 32,                           .data
		.lphy_avst_sink_dsp_capture_chan  (lphy_avst_sink_dsp_capture_channel),                               //   input,    width = 3,                           .channel
		.dxc_avst_sink_dsp_capture_valid  (dxc_avst_sink_dsp_capture_valid),                                  //   input,    width = 1,  dxc_avst_sink_dsp_capture.valid
		.dxc_avst_sink_dsp_capture_data   (dxc_avst_sink_dsp_capture_data),                                   //   input,   width = 32,                           .data
		.dxc_avst_sink_dsp_capture_chan   (dxc_avst_sink_dsp_capture_channel),                                //   input,    width = 3,                           .channel
		.interface_sel                    (interface_sel_data)                                                //  output,   width = 32,              interface_sel.data
	);

	ed_synth_clock_bridge_dsp clock_bridge_dsp (
		.in_clk  (dsp_in_clk_clk),               //   input,  width = 1,  in_clk.clk
		.out_clk (clock_bridge_dsp_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	ed_synth_clock_bridge_eth clock_bridge_eth (
		.in_clk  (eth_in_clk_clk),               //   input,  width = 1,  in_clk.clk
		.out_clk (clock_bridge_eth_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	clock_csr clock_csr (
		.in_clk  (clock_csr_clk),         //   input,  width = 1,  in_clk.clk
		.out_clk (clock_csr_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	ed_synth_clock_bridge_dspby2 ed_synth_clock_bridge_dspby2 (
		.in_clk  (clock_bridge_dspby2_in_clk_clk),           //   input,  width = 1,  in_clk.clk
		.out_clk (ed_synth_clock_bridge_dspby2_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	ed_synth_h2f_bridge ed_synth_h2f_bridge (
		.clk              (clock_csr_out_clk_clk),                //   input,    width = 1,   clk.clk
		.reset            (rst_controller_reset_out_reset),       //   input,    width = 1, reset.reset
		.s0_waitrequest   (ed_synth_h2f_bridge_s0_waitrequest),   //  output,    width = 1,    s0.waitrequest
		.s0_readdata      (ed_synth_h2f_bridge_s0_readdata),      //  output,  width = 512,      .readdata
		.s0_readdatavalid (ed_synth_h2f_bridge_s0_readdatavalid), //  output,    width = 1,      .readdatavalid
		.s0_burstcount    (ed_synth_h2f_bridge_s0_burstcount),    //   input,    width = 1,      .burstcount
		.s0_writedata     (ed_synth_h2f_bridge_s0_writedata),     //   input,  width = 512,      .writedata
		.s0_address       (ed_synth_h2f_bridge_s0_address),       //   input,   width = 28,      .address
		.s0_write         (ed_synth_h2f_bridge_s0_write),         //   input,    width = 1,      .write
		.s0_read          (ed_synth_h2f_bridge_s0_read),          //   input,    width = 1,      .read
		.s0_byteenable    (ed_synth_h2f_bridge_s0_byteenable),    //   input,   width = 64,      .byteenable
		.s0_debugaccess   (ed_synth_h2f_bridge_s0_debugaccess),   //   input,    width = 1,      .debugaccess
		.m0_waitrequest   (ed_synth_h2f_bridge_m0_waitrequest),   //   input,    width = 1,    m0.waitrequest
		.m0_readdata      (ed_synth_h2f_bridge_m0_readdata),      //   input,  width = 512,      .readdata
		.m0_readdatavalid (ed_synth_h2f_bridge_m0_readdatavalid), //   input,    width = 1,      .readdatavalid
		.m0_burstcount    (ed_synth_h2f_bridge_m0_burstcount),    //  output,    width = 1,      .burstcount
		.m0_writedata     (ed_synth_h2f_bridge_m0_writedata),     //  output,  width = 512,      .writedata
		.m0_address       (ed_synth_h2f_bridge_m0_address),       //  output,   width = 28,      .address
		.m0_write         (ed_synth_h2f_bridge_m0_write),         //  output,    width = 1,      .write
		.m0_read          (ed_synth_h2f_bridge_m0_read),          //  output,    width = 1,      .read
		.m0_byteenable    (ed_synth_h2f_bridge_m0_byteenable),    //  output,   width = 64,      .byteenable
		.m0_debugaccess   (ed_synth_h2f_bridge_m0_debugaccess)    //  output,    width = 1,      .debugaccess
	);

	ed_synth_h2f_lw_bridge ed_synth_h2f_lw_bridge (
		.clk              (clock_csr_out_clk_clk),                   //   input,   width = 1,   clk.clk
		.reset            (rst_controller_reset_out_reset),          //   input,   width = 1, reset.reset
		.s0_waitrequest   (h2f_lw_bridge_s0_waitrequest),            //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (h2f_lw_bridge_s0_readdata),               //  output,  width = 32,      .readdata
		.s0_readdatavalid (h2f_lw_bridge_s0_readdatavalid),          //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (h2f_lw_bridge_s0_burstcount),             //   input,   width = 1,      .burstcount
		.s0_writedata     (h2f_lw_bridge_s0_writedata),              //   input,  width = 32,      .writedata
		.s0_address       (h2f_lw_bridge_s0_address),                //   input,  width = 13,      .address
		.s0_write         (h2f_lw_bridge_s0_write),                  //   input,   width = 1,      .write
		.s0_read          (h2f_lw_bridge_s0_read),                   //   input,   width = 1,      .read
		.s0_byteenable    (h2f_lw_bridge_s0_byteenable),             //   input,   width = 4,      .byteenable
		.s0_debugaccess   (h2f_lw_bridge_s0_debugaccess),            //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (ed_synth_h2f_lw_bridge_m0_waitrequest),   //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (ed_synth_h2f_lw_bridge_m0_readdata),      //   input,  width = 32,      .readdata
		.m0_readdatavalid (ed_synth_h2f_lw_bridge_m0_readdatavalid), //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (ed_synth_h2f_lw_bridge_m0_burstcount),    //  output,   width = 1,      .burstcount
		.m0_writedata     (ed_synth_h2f_lw_bridge_m0_writedata),     //  output,  width = 32,      .writedata
		.m0_address       (ed_synth_h2f_lw_bridge_m0_address),       //  output,  width = 13,      .address
		.m0_write         (ed_synth_h2f_lw_bridge_m0_write),         //  output,   width = 1,      .write
		.m0_read          (ed_synth_h2f_lw_bridge_m0_read),          //  output,   width = 1,      .read
		.m0_byteenable    (ed_synth_h2f_lw_bridge_m0_byteenable),    //  output,   width = 4,      .byteenable
		.m0_debugaccess   (ed_synth_h2f_lw_bridge_m0_debugaccess)    //  output,   width = 1,      .debugaccess
	);

	ed_synth_reset_bridge_dsp ed_synth_reset_bridge_dsp (
		.clk         (clock_bridge_dsp_out_clk_clk),              //   input,  width = 1,       clk.clk
		.in_reset_n  (dsp_in_reset_reset_n),                      //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (ed_synth_reset_bridge_dsp_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	ed_synth_reset_bridge_eth ed_synth_reset_bridge_eth (
		.clk         (clock_bridge_eth_out_clk_clk),              //   input,  width = 1,       clk.clk
		.in_reset_n  (eth_in_reset_reset_n),                      //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (ed_synth_reset_bridge_eth_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	ed_synth_ninit_done_inst ninit_done_inst (
		.ninit_done ()  //  output,  width = 1, ninit_done.ninit_done
	);

	reset_csr reset_csr (
		.clk         (clock_csr_out_clk_clk),     //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_csr_reset_n),         //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (reset_csr_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	ddr4_wr_rd ddr4_wr_rd_0 (
		.emif_mm_slave_0_address        (),                                                             //   input,   width = 21,     emif_mm_slave_0.address
		.emif_mm_slave_0_read           (),                                                             //   input,    width = 1,                    .read
		.emif_mm_slave_0_readdata       (),                                                             //  output,  width = 128,                    .readdata
		.emif_mm_slave_0_write          (),                                                             //   input,    width = 1,                    .write
		.emif_mm_slave_0_writedata      (),                                                             //   input,  width = 128,                    .writedata
		.emif_mm_slave_0_readdatavalid  (),                                                             //  output,    width = 1,                    .readdatavalid
		.emif_mm_slave_0_waitrequest    (),                                                             //  output,    width = 1,                    .waitrequest
		.emif_mm_slave_0_byteenable     (),                                                             //   input,   width = 16,                    .byteenable
		.emif_mm_slave_0_burstcount     (),                                                             //   input,    width = 7,                    .burstcount
		.addr_span_0_cntl_read          (),                                                             //   input,    width = 1,    addr_span_0_cntl.read
		.addr_span_0_cntl_readdata      (),                                                             //  output,   width = 64,                    .readdata
		.addr_span_0_cntl_write         (),                                                             //   input,    width = 1,                    .write
		.addr_span_0_cntl_writedata     (),                                                             //   input,   width = 64,                    .writedata
		.addr_span_0_cntl_byteenable    (),                                                             //   input,    width = 8,                    .byteenable
		.emif_mm_slave_1_address        (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_address),       //   input,   width = 21,     emif_mm_slave_1.address
		.emif_mm_slave_1_read           (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_read),          //   input,    width = 1,                    .read
		.emif_mm_slave_1_readdata       (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_readdata),      //  output,  width = 128,                    .readdata
		.emif_mm_slave_1_write          (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_write),         //   input,    width = 1,                    .write
		.emif_mm_slave_1_writedata      (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_writedata),     //   input,  width = 128,                    .writedata
		.emif_mm_slave_1_readdatavalid  (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_readdatavalid), //  output,    width = 1,                    .readdatavalid
		.emif_mm_slave_1_waitrequest    (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_waitrequest),   //  output,    width = 1,                    .waitrequest
		.emif_mm_slave_1_byteenable     (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_byteenable),    //   input,   width = 16,                    .byteenable
		.emif_mm_slave_1_burstcount     (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_burstcount),    //   input,    width = 7,                    .burstcount
		.addr_span_1_cntl_read          (),                                                             //   input,    width = 1,    addr_span_1_cntl.read
		.addr_span_1_cntl_readdata      (),                                                             //  output,   width = 64,                    .readdata
		.addr_span_1_cntl_write         (),                                                             //   input,    width = 1,                    .write
		.addr_span_1_cntl_writedata     (),                                                             //   input,   width = 64,                    .writedata
		.addr_span_1_cntl_byteenable    (),                                                             //   input,    width = 8,                    .byteenable
		.wr_msgdma_ddr_address          (),                                                             //  output,   width = 32,       wr_msgdma_ddr.address
		.wr_msgdma_ddr_read             (),                                                             //  output,    width = 1,                    .read
		.wr_msgdma_ddr_waitrequest      (),                                                             //   input,    width = 1,                    .waitrequest
		.wr_msgdma_ddr_readdata         (),                                                             //   input,  width = 128,                    .readdata
		.wr_msgdma_ddr_write            (),                                                             //  output,    width = 1,                    .write
		.wr_msgdma_ddr_writedata        (),                                                             //  output,  width = 128,                    .writedata
		.wr_msgdma_ddr_readdatavalid    (),                                                             //   input,    width = 1,                    .readdatavalid
		.wr_msgdma_ddr_byteenable       (),                                                             //  output,   width = 16,                    .byteenable
		.wr_msgdma_ddr_burstcount       (),                                                             //  output,    width = 7,                    .burstcount
		.in_clk_clk                     (ed_synth_clock_bridge_dspby2_out_clk_clk),                     //   input,    width = 1,              in_clk.clk
		.csr_bridge_s0_waitrequest      (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_waitrequest),     //  output,    width = 1,       csr_bridge_s0.waitrequest
		.csr_bridge_s0_readdata         (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_readdata),        //  output,   width = 32,                    .readdata
		.csr_bridge_s0_readdatavalid    (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_readdatavalid),   //  output,    width = 1,                    .readdatavalid
		.csr_bridge_s0_burstcount       (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_burstcount),      //   input,    width = 1,                    .burstcount
		.csr_bridge_s0_writedata        (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_writedata),       //   input,   width = 32,                    .writedata
		.csr_bridge_s0_address          (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_address),         //   input,    width = 6,                    .address
		.csr_bridge_s0_write            (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_write),           //   input,    width = 1,                    .write
		.csr_bridge_s0_read             (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_read),            //   input,    width = 1,                    .read
		.csr_bridge_s0_byteenable       (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_byteenable),      //   input,    width = 4,                    .byteenable
		.csr_bridge_s0_debugaccess      (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_debugaccess),     //   input,    width = 1,                    .debugaccess
		.ocm_rd_address                 (mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_address),                //   input,   width = 13,              ocm_rd.address
		.ocm_rd_read                    (mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_read),                   //   input,    width = 1,                    .read
		.ocm_rd_readdata                (mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_readdata),               //  output,  width = 128,                    .readdata
		.ocm_rd_clk_clk                 (clock_csr_out_clk_clk),                                        //   input,    width = 1,          ocm_rd_clk.clk
		.ocm_rd_reset_reset             (rst_controller_reset_out_reset),                               //   input,    width = 1,        ocm_rd_reset.reset
		.ocm_rd_reset_reset_req         (rst_controller_reset_out_reset_req),                           //   input,    width = 1,                    .reset_req
		.emif_mm_master_1_waitrequest   (),                                                             //   input,    width = 1,    emif_mm_master_1.waitrequest
		.emif_mm_master_1_readdata      (),                                                             //   input,  width = 128,                    .readdata
		.emif_mm_master_1_readdatavalid (),                                                             //   input,    width = 1,                    .readdatavalid
		.emif_mm_master_1_burstcount    (),                                                             //  output,    width = 7,                    .burstcount
		.emif_mm_master_1_writedata     (),                                                             //  output,  width = 128,                    .writedata
		.emif_mm_master_1_address       (),                                                             //  output,   width = 10,                    .address
		.emif_mm_master_1_write         (),                                                             //  output,    width = 1,                    .write
		.emif_mm_master_1_read          (),                                                             //  output,    width = 1,                    .read
		.emif_mm_master_1_byteenable    (),                                                             //  output,   width = 16,                    .byteenable
		.emif_mm_master_1_debugaccess   (),                                                             //  output,    width = 1,                    .debugaccess
		.in_reset_reset_n               (~rst_controller_001_reset_out_reset),                          //   input,    width = 1,            in_reset.reset_n
		.wr_msgdma_0_csr_irq_irq        (wr_msgdma_0_csr_irq_irq),                                      //  output,    width = 1, wr_msgdma_0_csr_irq.irq
		.wr_msgdma_0_st_sink_data       (capture_if_top_0_avst_source_capture_data),                    //   input,  width = 128, wr_msgdma_0_st_sink.data
		.wr_msgdma_0_st_sink_valid      (capture_if_top_0_avst_source_capture_valid),                   //   input,    width = 1,                    .valid
		.wr_msgdma_0_st_sink_ready      (capture_if_top_0_avst_source_capture_ready)                    //  output,    width = 1,                    .ready
	);

	ed_synth_altera_mm_interconnect_1920_ff4yeri mm_interconnect_0 (
		.ed_synth_h2f_lw_bridge_m0_address                                       (ed_synth_h2f_lw_bridge_m0_address),                                //   input,  width = 13,                                         ed_synth_h2f_lw_bridge_m0.address
		.ed_synth_h2f_lw_bridge_m0_waitrequest                                   (ed_synth_h2f_lw_bridge_m0_waitrequest),                            //  output,   width = 1,                                                                  .waitrequest
		.ed_synth_h2f_lw_bridge_m0_burstcount                                    (ed_synth_h2f_lw_bridge_m0_burstcount),                             //   input,   width = 1,                                                                  .burstcount
		.ed_synth_h2f_lw_bridge_m0_byteenable                                    (ed_synth_h2f_lw_bridge_m0_byteenable),                             //   input,   width = 4,                                                                  .byteenable
		.ed_synth_h2f_lw_bridge_m0_read                                          (ed_synth_h2f_lw_bridge_m0_read),                                   //   input,   width = 1,                                                                  .read
		.ed_synth_h2f_lw_bridge_m0_readdata                                      (ed_synth_h2f_lw_bridge_m0_readdata),                               //  output,  width = 32,                                                                  .readdata
		.ed_synth_h2f_lw_bridge_m0_readdatavalid                                 (ed_synth_h2f_lw_bridge_m0_readdatavalid),                          //  output,   width = 1,                                                                  .readdatavalid
		.ed_synth_h2f_lw_bridge_m0_write                                         (ed_synth_h2f_lw_bridge_m0_write),                                  //   input,   width = 1,                                                                  .write
		.ed_synth_h2f_lw_bridge_m0_writedata                                     (ed_synth_h2f_lw_bridge_m0_writedata),                              //   input,  width = 32,                                                                  .writedata
		.ed_synth_h2f_lw_bridge_m0_debugaccess                                   (ed_synth_h2f_lw_bridge_m0_debugaccess),                            //   input,   width = 1,                                                                  .debugaccess
		.ddr4_wr_rd_0_csr_bridge_s0_address                                      (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_address),             //  output,   width = 6,                                        ddr4_wr_rd_0_csr_bridge_s0.address
		.ddr4_wr_rd_0_csr_bridge_s0_write                                        (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_write),               //  output,   width = 1,                                                                  .write
		.ddr4_wr_rd_0_csr_bridge_s0_read                                         (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_read),                //  output,   width = 1,                                                                  .read
		.ddr4_wr_rd_0_csr_bridge_s0_readdata                                     (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_readdata),            //   input,  width = 32,                                                                  .readdata
		.ddr4_wr_rd_0_csr_bridge_s0_writedata                                    (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_writedata),           //  output,  width = 32,                                                                  .writedata
		.ddr4_wr_rd_0_csr_bridge_s0_burstcount                                   (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_burstcount),          //  output,   width = 1,                                                                  .burstcount
		.ddr4_wr_rd_0_csr_bridge_s0_byteenable                                   (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_byteenable),          //  output,   width = 4,                                                                  .byteenable
		.ddr4_wr_rd_0_csr_bridge_s0_readdatavalid                                (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_readdatavalid),       //   input,   width = 1,                                                                  .readdatavalid
		.ddr4_wr_rd_0_csr_bridge_s0_waitrequest                                  (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_waitrequest),         //   input,   width = 1,                                                                  .waitrequest
		.ddr4_wr_rd_0_csr_bridge_s0_debugaccess                                  (mm_interconnect_0_ddr4_wr_rd_0_csr_bridge_s0_debugaccess),         //  output,   width = 1,                                                                  .debugaccess
		.capture_if_top_0_csr_dsp_capture_address                                (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_address),       //  output,   width = 5,                                  capture_if_top_0_csr_dsp_capture.address
		.capture_if_top_0_csr_dsp_capture_write                                  (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_write),         //  output,   width = 1,                                                                  .write
		.capture_if_top_0_csr_dsp_capture_read                                   (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_read),          //  output,   width = 1,                                                                  .read
		.capture_if_top_0_csr_dsp_capture_readdata                               (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_readdata),      //   input,  width = 32,                                                                  .readdata
		.capture_if_top_0_csr_dsp_capture_writedata                              (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_writedata),     //  output,  width = 32,                                                                  .writedata
		.capture_if_top_0_csr_dsp_capture_readdatavalid                          (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_readdatavalid), //   input,   width = 1,                                                                  .readdatavalid
		.capture_if_top_0_csr_dsp_capture_waitrequest                            (mm_interconnect_0_capture_if_top_0_csr_dsp_capture_waitrequest),   //   input,   width = 1,                                                                  .waitrequest
		.ed_synth_h2f_lw_bridge_reset_reset_bridge_in_reset_reset                (rst_controller_002_reset_out_reset),                               //   input,   width = 1,                ed_synth_h2f_lw_bridge_reset_reset_bridge_in_reset.reset
		.ddr4_wr_rd_0_in_reset_reset_bridge_in_reset_reset                       (rst_controller_003_reset_out_reset),                               //   input,   width = 1,                       ddr4_wr_rd_0_in_reset_reset_bridge_in_reset.reset
		.ed_synth_h2f_lw_bridge_m0_translator_reset_reset_bridge_in_reset_reset  (rst_controller_002_reset_out_reset),                               //   input,   width = 1,  ed_synth_h2f_lw_bridge_m0_translator_reset_reset_bridge_in_reset.reset
		.ddr4_wr_rd_0_csr_bridge_s0_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                               //   input,   width = 1, ddr4_wr_rd_0_csr_bridge_s0_translator_reset_reset_bridge_in_reset.reset
		.clock_csr_out_clk_clk                                                   (clock_csr_out_clk_clk),                                            //   input,   width = 1,                                                 clock_csr_out_clk.clk
		.ed_synth_clock_bridge_dspby2_out_clk_clk                                (ed_synth_clock_bridge_dspby2_out_clk_clk)                          //   input,   width = 1,                              ed_synth_clock_bridge_dspby2_out_clk.clk
	);

	ed_synth_altera_mm_interconnect_1920_urzwi2q mm_interconnect_1 (
		.ed_synth_h2f_bridge_m0_address                                            (ed_synth_h2f_bridge_m0_address),                               //   input,   width = 28,                                              ed_synth_h2f_bridge_m0.address
		.ed_synth_h2f_bridge_m0_waitrequest                                        (ed_synth_h2f_bridge_m0_waitrequest),                           //  output,    width = 1,                                                                    .waitrequest
		.ed_synth_h2f_bridge_m0_burstcount                                         (ed_synth_h2f_bridge_m0_burstcount),                            //   input,    width = 1,                                                                    .burstcount
		.ed_synth_h2f_bridge_m0_byteenable                                         (ed_synth_h2f_bridge_m0_byteenable),                            //   input,   width = 64,                                                                    .byteenable
		.ed_synth_h2f_bridge_m0_read                                               (ed_synth_h2f_bridge_m0_read),                                  //   input,    width = 1,                                                                    .read
		.ed_synth_h2f_bridge_m0_readdata                                           (ed_synth_h2f_bridge_m0_readdata),                              //  output,  width = 512,                                                                    .readdata
		.ed_synth_h2f_bridge_m0_readdatavalid                                      (ed_synth_h2f_bridge_m0_readdatavalid),                         //  output,    width = 1,                                                                    .readdatavalid
		.ed_synth_h2f_bridge_m0_write                                              (ed_synth_h2f_bridge_m0_write),                                 //   input,    width = 1,                                                                    .write
		.ed_synth_h2f_bridge_m0_writedata                                          (ed_synth_h2f_bridge_m0_writedata),                             //   input,  width = 512,                                                                    .writedata
		.ed_synth_h2f_bridge_m0_debugaccess                                        (ed_synth_h2f_bridge_m0_debugaccess),                           //   input,    width = 1,                                                                    .debugaccess
		.ddr4_wr_rd_0_emif_mm_slave_1_address                                      (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_address),       //  output,   width = 21,                                        ddr4_wr_rd_0_emif_mm_slave_1.address
		.ddr4_wr_rd_0_emif_mm_slave_1_write                                        (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_write),         //  output,    width = 1,                                                                    .write
		.ddr4_wr_rd_0_emif_mm_slave_1_read                                         (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_read),          //  output,    width = 1,                                                                    .read
		.ddr4_wr_rd_0_emif_mm_slave_1_readdata                                     (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_readdata),      //   input,  width = 128,                                                                    .readdata
		.ddr4_wr_rd_0_emif_mm_slave_1_writedata                                    (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_writedata),     //  output,  width = 128,                                                                    .writedata
		.ddr4_wr_rd_0_emif_mm_slave_1_burstcount                                   (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_burstcount),    //  output,    width = 7,                                                                    .burstcount
		.ddr4_wr_rd_0_emif_mm_slave_1_byteenable                                   (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_byteenable),    //  output,   width = 16,                                                                    .byteenable
		.ddr4_wr_rd_0_emif_mm_slave_1_readdatavalid                                (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_readdatavalid), //   input,    width = 1,                                                                    .readdatavalid
		.ddr4_wr_rd_0_emif_mm_slave_1_waitrequest                                  (mm_interconnect_1_ddr4_wr_rd_0_emif_mm_slave_1_waitrequest),   //   input,    width = 1,                                                                    .waitrequest
		.ddr4_wr_rd_0_ocm_rd_address                                               (mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_address),                //  output,   width = 13,                                                 ddr4_wr_rd_0_ocm_rd.address
		.ddr4_wr_rd_0_ocm_rd_read                                                  (mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_read),                   //  output,    width = 1,                                                                    .read
		.ddr4_wr_rd_0_ocm_rd_readdata                                              (mm_interconnect_1_ddr4_wr_rd_0_ocm_rd_readdata),               //   input,  width = 128,                                                                    .readdata
		.ed_synth_h2f_bridge_reset_reset_bridge_in_reset_reset                     (rst_controller_002_reset_out_reset),                           //   input,    width = 1,                     ed_synth_h2f_bridge_reset_reset_bridge_in_reset.reset
		.ddr4_wr_rd_0_in_reset_reset_bridge_in_reset_reset                         (rst_controller_003_reset_out_reset),                           //   input,    width = 1,                         ddr4_wr_rd_0_in_reset_reset_bridge_in_reset.reset
		.ed_synth_h2f_bridge_m0_translator_reset_reset_bridge_in_reset_reset       (rst_controller_002_reset_out_reset),                           //   input,    width = 1,       ed_synth_h2f_bridge_m0_translator_reset_reset_bridge_in_reset.reset
		.ddr4_wr_rd_0_emif_mm_slave_1_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                           //   input,    width = 1, ddr4_wr_rd_0_emif_mm_slave_1_translator_reset_reset_bridge_in_reset.reset
		.clock_csr_out_clk_clk                                                     (clock_csr_out_clk_clk),                                        //   input,    width = 1,                                                   clock_csr_out_clk.clk
		.ed_synth_clock_bridge_dspby2_out_clk_clk                                  (ed_synth_clock_bridge_dspby2_out_clk_clk)                      //   input,    width = 1,                                ed_synth_clock_bridge_dspby2_out_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_csr_out_reset_reset),         //   input,  width = 1, reset_in0.reset
		.clk            (clock_csr_out_clk_clk),              //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_csr_out_reset_reset),               //   input,  width = 1, reset_in0.reset
		.clk            (ed_synth_clock_bridge_dspby2_out_clk_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),       //  output,  width = 1, reset_out.reset
		.reset_req      (),                                         // (terminated),                       
		.reset_req_in0  (1'b0),                                     // (terminated),                       
		.reset_in1      (1'b0),                                     // (terminated),                       
		.reset_req_in1  (1'b0),                                     // (terminated),                       
		.reset_in2      (1'b0),                                     // (terminated),                       
		.reset_req_in2  (1'b0),                                     // (terminated),                       
		.reset_in3      (1'b0),                                     // (terminated),                       
		.reset_req_in3  (1'b0),                                     // (terminated),                       
		.reset_in4      (1'b0),                                     // (terminated),                       
		.reset_req_in4  (1'b0),                                     // (terminated),                       
		.reset_in5      (1'b0),                                     // (terminated),                       
		.reset_req_in5  (1'b0),                                     // (terminated),                       
		.reset_in6      (1'b0),                                     // (terminated),                       
		.reset_req_in6  (1'b0),                                     // (terminated),                       
		.reset_in7      (1'b0),                                     // (terminated),                       
		.reset_req_in7  (1'b0),                                     // (terminated),                       
		.reset_in8      (1'b0),                                     // (terminated),                       
		.reset_req_in8  (1'b0),                                     // (terminated),                       
		.reset_in9      (1'b0),                                     // (terminated),                       
		.reset_req_in9  (1'b0),                                     // (terminated),                       
		.reset_in10     (1'b0),                                     // (terminated),                       
		.reset_req_in10 (1'b0),                                     // (terminated),                       
		.reset_in11     (1'b0),                                     // (terminated),                       
		.reset_req_in11 (1'b0),                                     // (terminated),                       
		.reset_in12     (1'b0),                                     // (terminated),                       
		.reset_req_in12 (1'b0),                                     // (terminated),                       
		.reset_in13     (1'b0),                                     // (terminated),                       
		.reset_req_in13 (1'b0),                                     // (terminated),                       
		.reset_in14     (1'b0),                                     // (terminated),                       
		.reset_req_in14 (1'b0),                                     // (terminated),                       
		.reset_in15     (1'b0),                                     // (terminated),                       
		.reset_req_in15 (1'b0)                                      // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_csr_out_reset_reset),         //   input,  width = 1, reset_in0.reset
		.clk            (clock_csr_out_clk_clk),              //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_csr_out_reset_reset),               //   input,  width = 1, reset_in0.reset
		.clk            (ed_synth_clock_bridge_dspby2_out_clk_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),       //  output,  width = 1, reset_out.reset
		.reset_req      (),                                         // (terminated),                       
		.reset_req_in0  (1'b0),                                     // (terminated),                       
		.reset_in1      (1'b0),                                     // (terminated),                       
		.reset_req_in1  (1'b0),                                     // (terminated),                       
		.reset_in2      (1'b0),                                     // (terminated),                       
		.reset_req_in2  (1'b0),                                     // (terminated),                       
		.reset_in3      (1'b0),                                     // (terminated),                       
		.reset_req_in3  (1'b0),                                     // (terminated),                       
		.reset_in4      (1'b0),                                     // (terminated),                       
		.reset_req_in4  (1'b0),                                     // (terminated),                       
		.reset_in5      (1'b0),                                     // (terminated),                       
		.reset_req_in5  (1'b0),                                     // (terminated),                       
		.reset_in6      (1'b0),                                     // (terminated),                       
		.reset_req_in6  (1'b0),                                     // (terminated),                       
		.reset_in7      (1'b0),                                     // (terminated),                       
		.reset_req_in7  (1'b0),                                     // (terminated),                       
		.reset_in8      (1'b0),                                     // (terminated),                       
		.reset_req_in8  (1'b0),                                     // (terminated),                       
		.reset_in9      (1'b0),                                     // (terminated),                       
		.reset_req_in9  (1'b0),                                     // (terminated),                       
		.reset_in10     (1'b0),                                     // (terminated),                       
		.reset_req_in10 (1'b0),                                     // (terminated),                       
		.reset_in11     (1'b0),                                     // (terminated),                       
		.reset_req_in11 (1'b0),                                     // (terminated),                       
		.reset_in12     (1'b0),                                     // (terminated),                       
		.reset_req_in12 (1'b0),                                     // (terminated),                       
		.reset_in13     (1'b0),                                     // (terminated),                       
		.reset_req_in13 (1'b0),                                     // (terminated),                       
		.reset_in14     (1'b0),                                     // (terminated),                       
		.reset_req_in14 (1'b0),                                     // (terminated),                       
		.reset_in15     (1'b0),                                     // (terminated),                       
		.reset_req_in15 (1'b0)                                      // (terminated),                       
	);

endmodule
