//`define SCH_LOOPBACK
//`define IFFT_FFT_LOOPBACK
//`define SHORT_PRACH_FORMAT
//`define OCM_CAPTURE
//`define CONFIG_CC1
//`define CONFIG_CC2
