// subsys_ftile_25gbe_1588.v

// Generated using ACDS version 24.1 115

`timescale 1 ps / 1 ps
module subsys_ftile_25gbe_1588 #(
		parameter FP_WIDTH = 8
	) (
		input  wire         rx_dma_resetn,                                               //                                   rx_dma_resetn.reset_n
		output wire         csr_waitrequest,                                             //                                             csr.waitrequest
		output wire [31:0]  csr_readdata,                                                //                                                .readdata
		output wire         csr_readdatavalid,                                           //                                                .readdatavalid
		input  wire [0:0]   csr_burstcount,                                              //                                                .burstcount
		input  wire [31:0]  csr_writedata,                                               //                                                .writedata
		input  wire [7:0]   csr_address,                                                 //                                                .address
		input  wire         csr_write,                                                   //                                                .write
		input  wire         csr_read,                                                    //                                                .read
		input  wire [3:0]   csr_byteenable,                                              //                                                .byteenable
		input  wire         csr_debugaccess,                                             //                                                .debugaccess
		input  wire         clk_clk,                                                     //                                             clk.clk
		input  wire         subsys_ftile_25gbe_1588_dmaclkout_in_clk_clk,                //        subsys_ftile_25gbe_1588_dmaclkout_in_clk.clk
		input  wire         subsys_ftile_25gbe_1588_o_pll_clk_in_clk_clk,                //        subsys_ftile_25gbe_1588_o_pll_clk_in_clk.clk
		input  wire         reset_reset_n,                                               //                                           reset.reset_n
		input  wire         ftile_25gbe_rx_dma_ch1_pktin_startofpacket,                  //                    ftile_25gbe_rx_dma_ch1_pktin.startofpacket
		input  wire         ftile_25gbe_rx_dma_ch1_pktin_valid,                          //                                                .valid
		input  wire         ftile_25gbe_rx_dma_ch1_pktin_endofpacket,                    //                                                .endofpacket
		input  wire [63:0]  ftile_25gbe_rx_dma_ch1_pktin_data,                           //                                                .data
		input  wire [2:0]   ftile_25gbe_rx_dma_ch1_pktin_empty,                          //                                                .empty
		input  wire [5:0]   ftile_25gbe_rx_dma_ch1_pktin_error,                          //                                                .error
		input  wire         ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_valid,            //      ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts.valid
		input  wire [95:0]  ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_data,             //                                                .data
		output wire [36:0]  rx_dma_ch1_prefetcher_read_master_address,                   //               rx_dma_ch1_prefetcher_read_master.address
		output wire         rx_dma_ch1_prefetcher_read_master_read,                      //                                                .read
		input  wire [127:0] rx_dma_ch1_prefetcher_read_master_readdata,                  //                                                .readdata
		input  wire         rx_dma_ch1_prefetcher_read_master_waitrequest,               //                                                .waitrequest
		input  wire         rx_dma_ch1_prefetcher_read_master_readdatavalid,             //                                                .readdatavalid
		output wire [2:0]   rx_dma_ch1_prefetcher_read_master_burstcount,                //                                                .burstcount
		output wire [36:0]  rx_dma_ch1_prefetcher_write_master_address,                  //              rx_dma_ch1_prefetcher_write_master.address
		output wire         rx_dma_ch1_prefetcher_write_master_write,                    //                                                .write
		output wire [15:0]  rx_dma_ch1_prefetcher_write_master_byteenable,               //                                                .byteenable
		output wire [127:0] rx_dma_ch1_prefetcher_write_master_writedata,                //                                                .writedata
		input  wire         rx_dma_ch1_prefetcher_write_master_waitrequest,              //                                                .waitrequest
		input  wire [1:0]   rx_dma_ch1_prefetcher_write_master_response,                 //                                                .response
		input  wire         rx_dma_ch1_prefetcher_write_master_writeresponsevalid,       //                                                .writeresponsevalid
		output wire         rx_dma_ch1_irq_irq,                                          //                                  rx_dma_ch1_irq.irq
		output wire [36:0]  rx_dma_ch1_write_master_address,                             //                         rx_dma_ch1_write_master.address
		output wire         rx_dma_ch1_write_master_write,                               //                                                .write
		output wire [15:0]  rx_dma_ch1_write_master_byteenable,                          //                                                .byteenable
		output wire [127:0] rx_dma_ch1_write_master_writedata,                           //                                                .writedata
		input  wire         rx_dma_ch1_write_master_waitrequest,                         //                                                .waitrequest
		output wire [4:0]   rx_dma_ch1_write_master_burstcount,                          //                                                .burstcount
		input  wire [1:0]   rx_dma_ch1_write_master_response,                            //                                                .response
		input  wire         rx_dma_ch1_write_master_writeresponsevalid,                  //                                                .writeresponsevalid
		input  wire [0:0]   ts_chs_compl_0_clk_bus_in_clk,                               //                       ts_chs_compl_0_clk_bus_in.clk
		input  wire [0:0]   ts_chs_compl_0_rst_bus_in_reset,                             //                       ts_chs_compl_0_rst_bus_in.reset
		input  wire [0:0]   ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_valid,            //      ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts.valid
		input  wire [19:0]  ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_fingerprint,      //                                                .fingerprint
		input  wire [95:0]  ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_data,             //                                                .data
		input  wire         ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready,           //     ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st.ready
		output wire         ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket,   //                                                .startofpacket
		output wire         ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid,           //                                                .valid
		output wire         ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket,     //                                                .endofpacket
		output wire [63:0]  ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data,            //                                                .data
		output wire [2:0]   ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty,           //                                                .empty
		output wire [0:0]   ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error,           //                                                .error
		output wire         ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_valid,       // ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req.valid
		output wire [19:0]  ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_fingerprint, //                                                .fingerprint
		output wire [36:0]  tx_dma_ch1_prefetcher_read_master_address,                   //               tx_dma_ch1_prefetcher_read_master.address
		output wire         tx_dma_ch1_prefetcher_read_master_read,                      //                                                .read
		input  wire [127:0] tx_dma_ch1_prefetcher_read_master_readdata,                  //                                                .readdata
		input  wire         tx_dma_ch1_prefetcher_read_master_waitrequest,               //                                                .waitrequest
		input  wire         tx_dma_ch1_prefetcher_read_master_readdatavalid,             //                                                .readdatavalid
		output wire [2:0]   tx_dma_ch1_prefetcher_read_master_burstcount,                //                                                .burstcount
		output wire [36:0]  tx_dma_ch1_prefetcher_write_master_address,                  //              tx_dma_ch1_prefetcher_write_master.address
		output wire         tx_dma_ch1_prefetcher_write_master_write,                    //                                                .write
		output wire [15:0]  tx_dma_ch1_prefetcher_write_master_byteenable,               //                                                .byteenable
		output wire [127:0] tx_dma_ch1_prefetcher_write_master_writedata,                //                                                .writedata
		input  wire         tx_dma_ch1_prefetcher_write_master_waitrequest,              //                                                .waitrequest
		input  wire [1:0]   tx_dma_ch1_prefetcher_write_master_response,                 //                                                .response
		input  wire         tx_dma_ch1_prefetcher_write_master_writeresponsevalid,       //                                                .writeresponsevalid
		output wire         tx_dma_ch1_irq_irq,                                          //                                  tx_dma_ch1_irq.irq
		output wire [36:0]  tx_dma_ch1_read_master_address,                              //                          tx_dma_ch1_read_master.address
		output wire         tx_dma_ch1_read_master_read,                                 //                                                .read
		output wire [15:0]  tx_dma_ch1_read_master_byteenable,                           //                                                .byteenable
		input  wire [127:0] tx_dma_ch1_read_master_readdata,                             //                                                .readdata
		input  wire         tx_dma_ch1_read_master_waitrequest,                          //                                                .waitrequest
		input  wire         tx_dma_ch1_read_master_readdatavalid,                        //                                                .readdatavalid
		output wire [4:0]   tx_dma_ch1_read_master_burstcount                            //                                                .burstcount
	);

	wire         subsys_ftile_25gbe_1588_csrclk_out_clk_clk;                 // subsys_ftile_25gbe_1588_csrclk:out_clk -> [mm_interconnect_0:subsys_ftile_25gbe_1588_csrclk_out_clk_clk, subsys_ftile_25gbe_1588_csr:clk, subsys_ftile_25gbe_1588_reset:clk]
	wire         subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk;              // subsys_ftile_25gbe_1588_dmaclkout:out_clk -> [ftile_25gbe_rx_dma_ch1:dma_clk_clk, ftile_25gbe_tx_dma_ch1:dma_clk_clk, mm_interconnect_0:subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk, rst_controller:clk, rx_dma_reset_bridge:clk]
	wire         subsys_ftile_25gbe_1588_o_pll_clk_out_clk_clk;              // subsys_ftile_25gbe_1588_o_pll_clk:out_clk -> [ftile_25gbe_rx_dma_ch1:ftile_clk_clk, ftile_25gbe_tx_dma_ch1:ftile_clk_clk]
	wire         subsys_ftile_25gbe_1588_reset_out_reset_reset;              // subsys_ftile_25gbe_1588_reset:out_reset_n -> [mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:subsys_ftile_25gbe_1588_csr_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0, subsys_ftile_25gbe_1588_csr:reset]
	wire         rx_dma_reset_bridge_out_reset_reset;                        // rx_dma_reset_bridge:out_reset_n -> [ftile_25gbe_rx_dma_ch1:reset_reset_n, mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_agent_rsp_fifo_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:ftile_25gbe_rx_dma_ch1_reset_reset_bridge_in_reset_reset]
	wire         subsys_ftile_25gbe_1588_csr_m0_waitrequest;                 // mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_waitrequest -> subsys_ftile_25gbe_1588_csr:m0_waitrequest
	wire  [31:0] subsys_ftile_25gbe_1588_csr_m0_readdata;                    // mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_readdata -> subsys_ftile_25gbe_1588_csr:m0_readdata
	wire         subsys_ftile_25gbe_1588_csr_m0_debugaccess;                 // subsys_ftile_25gbe_1588_csr:m0_debugaccess -> mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_debugaccess
	wire   [7:0] subsys_ftile_25gbe_1588_csr_m0_address;                     // subsys_ftile_25gbe_1588_csr:m0_address -> mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_address
	wire         subsys_ftile_25gbe_1588_csr_m0_read;                        // subsys_ftile_25gbe_1588_csr:m0_read -> mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_read
	wire   [3:0] subsys_ftile_25gbe_1588_csr_m0_byteenable;                  // subsys_ftile_25gbe_1588_csr:m0_byteenable -> mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_byteenable
	wire         subsys_ftile_25gbe_1588_csr_m0_readdatavalid;               // mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_readdatavalid -> subsys_ftile_25gbe_1588_csr:m0_readdatavalid
	wire  [31:0] subsys_ftile_25gbe_1588_csr_m0_writedata;                   // subsys_ftile_25gbe_1588_csr:m0_writedata -> mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_writedata
	wire         subsys_ftile_25gbe_1588_csr_m0_write;                       // subsys_ftile_25gbe_1588_csr:m0_write -> mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_write
	wire   [0:0] subsys_ftile_25gbe_1588_csr_m0_burstcount;                  // subsys_ftile_25gbe_1588_csr:m0_burstcount -> mm_interconnect_0:subsys_ftile_25gbe_1588_csr_m0_burstcount
	wire  [31:0] mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_readdata;      // ftile_25gbe_tx_dma_ch1:csr_readdata -> mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_readdata
	wire         mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_waitrequest;   // ftile_25gbe_tx_dma_ch1:csr_waitrequest -> mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_waitrequest
	wire         mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_debugaccess;   // mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_debugaccess -> ftile_25gbe_tx_dma_ch1:csr_debugaccess
	wire   [5:0] mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_address;       // mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_address -> ftile_25gbe_tx_dma_ch1:csr_address
	wire         mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_read;          // mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_read -> ftile_25gbe_tx_dma_ch1:csr_read
	wire   [3:0] mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_byteenable;    // mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_byteenable -> ftile_25gbe_tx_dma_ch1:csr_byteenable
	wire         mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_readdatavalid; // ftile_25gbe_tx_dma_ch1:csr_readdatavalid -> mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_readdatavalid
	wire         mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_write;         // mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_write -> ftile_25gbe_tx_dma_ch1:csr_write
	wire  [31:0] mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_writedata;     // mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_writedata -> ftile_25gbe_tx_dma_ch1:csr_writedata
	wire   [0:0] mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_burstcount;    // mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_burstcount -> ftile_25gbe_tx_dma_ch1:csr_burstcount
	wire  [31:0] mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_readdata;      // ftile_25gbe_rx_dma_ch1:csr_readdata -> mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_readdata
	wire         mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_waitrequest;   // ftile_25gbe_rx_dma_ch1:csr_waitrequest -> mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_waitrequest
	wire         mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_debugaccess;   // mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_debugaccess -> ftile_25gbe_rx_dma_ch1:csr_debugaccess
	wire   [5:0] mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_address;       // mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_address -> ftile_25gbe_rx_dma_ch1:csr_address
	wire         mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_read;          // mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_read -> ftile_25gbe_rx_dma_ch1:csr_read
	wire   [3:0] mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_byteenable;    // mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_byteenable -> ftile_25gbe_rx_dma_ch1:csr_byteenable
	wire         mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_readdatavalid; // ftile_25gbe_rx_dma_ch1:csr_readdatavalid -> mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_readdatavalid
	wire         mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_write;         // mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_write -> ftile_25gbe_rx_dma_ch1:csr_write
	wire  [31:0] mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_writedata;     // mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_writedata -> ftile_25gbe_rx_dma_ch1:csr_writedata
	wire   [0:0] mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_burstcount;    // mm_interconnect_0:ftile_25gbe_rx_dma_ch1_csr_burstcount -> ftile_25gbe_rx_dma_ch1:csr_burstcount
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [ftile_25gbe_tx_dma_ch1:reset_reset_n, mm_interconnect_0:ftile_25gbe_tx_dma_ch1_csr_agent_rsp_fifo_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:ftile_25gbe_tx_dma_ch1_reset_reset_bridge_in_reset_reset]

	rx_dma_reset_bridge rx_dma_reset_bridge (
		.clk         (subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk), //   input,  width = 1,       clk.clk
		.in_reset_n  (rx_dma_resetn),                                 //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (rx_dma_reset_bridge_out_reset_reset)            //  output,  width = 1, out_reset.reset_n
	);

	subsys_ftile_25gbe_1588_csr subsys_ftile_25gbe_1588_csr (
		.clk              (subsys_ftile_25gbe_1588_csrclk_out_clk_clk),     //   input,   width = 1,   clk.clk
		.reset            (~subsys_ftile_25gbe_1588_reset_out_reset_reset), //   input,   width = 1, reset.reset
		.s0_waitrequest   (csr_waitrequest),                                //  output,   width = 1,    s0.waitrequest
		.s0_readdata      (csr_readdata),                                   //  output,  width = 32,      .readdata
		.s0_readdatavalid (csr_readdatavalid),                              //  output,   width = 1,      .readdatavalid
		.s0_burstcount    (csr_burstcount),                                 //   input,   width = 1,      .burstcount
		.s0_writedata     (csr_writedata),                                  //   input,  width = 32,      .writedata
		.s0_address       (csr_address),                                    //   input,   width = 8,      .address
		.s0_write         (csr_write),                                      //   input,   width = 1,      .write
		.s0_read          (csr_read),                                       //   input,   width = 1,      .read
		.s0_byteenable    (csr_byteenable),                                 //   input,   width = 4,      .byteenable
		.s0_debugaccess   (csr_debugaccess),                                //   input,   width = 1,      .debugaccess
		.m0_waitrequest   (subsys_ftile_25gbe_1588_csr_m0_waitrequest),     //   input,   width = 1,    m0.waitrequest
		.m0_readdata      (subsys_ftile_25gbe_1588_csr_m0_readdata),        //   input,  width = 32,      .readdata
		.m0_readdatavalid (subsys_ftile_25gbe_1588_csr_m0_readdatavalid),   //   input,   width = 1,      .readdatavalid
		.m0_burstcount    (subsys_ftile_25gbe_1588_csr_m0_burstcount),      //  output,   width = 1,      .burstcount
		.m0_writedata     (subsys_ftile_25gbe_1588_csr_m0_writedata),       //  output,  width = 32,      .writedata
		.m0_address       (subsys_ftile_25gbe_1588_csr_m0_address),         //  output,   width = 8,      .address
		.m0_write         (subsys_ftile_25gbe_1588_csr_m0_write),           //  output,   width = 1,      .write
		.m0_read          (subsys_ftile_25gbe_1588_csr_m0_read),            //  output,   width = 1,      .read
		.m0_byteenable    (subsys_ftile_25gbe_1588_csr_m0_byteenable),      //  output,   width = 4,      .byteenable
		.m0_debugaccess   (subsys_ftile_25gbe_1588_csr_m0_debugaccess)      //  output,   width = 1,      .debugaccess
	);

	subsys_ftile_25gbe_1588_csrclk subsys_ftile_25gbe_1588_csrclk (
		.in_clk  (clk_clk),                                    //   input,  width = 1,  in_clk.clk
		.out_clk (subsys_ftile_25gbe_1588_csrclk_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	subsys_ftile_25gbe_1588_dmaclkout subsys_ftile_25gbe_1588_dmaclkout (
		.in_clk  (subsys_ftile_25gbe_1588_dmaclkout_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	subsys_ftile_25gbe_1588_o_pll_clk subsys_ftile_25gbe_1588_o_pll_clk (
		.in_clk  (subsys_ftile_25gbe_1588_o_pll_clk_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (subsys_ftile_25gbe_1588_o_pll_clk_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	subsys_ftile_25gbe_1588_reset subsys_ftile_25gbe_1588_reset (
		.clk         (subsys_ftile_25gbe_1588_csrclk_out_clk_clk),    //   input,  width = 1,       clk.clk
		.in_reset_n  (reset_reset_n),                                 //   input,  width = 1,  in_reset.reset_n
		.out_reset_n (subsys_ftile_25gbe_1588_reset_out_reset_reset)  //  output,  width = 1, out_reset.reset_n
	);

	subsys_ftile_25gbe_rx_dma ftile_25gbe_rx_dma_ch1 (
		.dma_clk_clk                                (subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk),              //   input,    width = 1,                 dma_clk.clk
		.csr_waitrequest                            (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_waitrequest),   //  output,    width = 1,                     csr.waitrequest
		.csr_readdata                               (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_readdata),      //  output,   width = 32,                        .readdata
		.csr_readdatavalid                          (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_readdatavalid), //  output,    width = 1,                        .readdatavalid
		.csr_burstcount                             (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_burstcount),    //   input,    width = 1,                        .burstcount
		.csr_writedata                              (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_writedata),     //   input,   width = 32,                        .writedata
		.csr_address                                (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_address),       //   input,    width = 6,                        .address
		.csr_write                                  (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_write),         //   input,    width = 1,                        .write
		.csr_read                                   (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_read),          //   input,    width = 1,                        .read
		.csr_byteenable                             (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_byteenable),    //   input,    width = 4,                        .byteenable
		.csr_debugaccess                            (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_debugaccess),   //   input,    width = 1,                        .debugaccess
		.pktin_startofpacket                        (ftile_25gbe_rx_dma_ch1_pktin_startofpacket),                 //   input,    width = 1,                   pktin.startofpacket
		.pktin_valid                                (ftile_25gbe_rx_dma_ch1_pktin_valid),                         //   input,    width = 1,                        .valid
		.pktin_endofpacket                          (ftile_25gbe_rx_dma_ch1_pktin_endofpacket),                   //   input,    width = 1,                        .endofpacket
		.pktin_data                                 (ftile_25gbe_rx_dma_ch1_pktin_data),                          //   input,   width = 64,                        .data
		.pktin_empty                                (ftile_25gbe_rx_dma_ch1_pktin_empty),                         //   input,    width = 3,                        .empty
		.pktin_error                                (ftile_25gbe_rx_dma_ch1_pktin_error),                         //   input,    width = 6,                        .error
		.rx_dma_fifo_0_in_ts_valid                  (ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_valid),           //   input,    width = 1,     rx_dma_fifo_0_in_ts.valid
		.rx_dma_fifo_0_in_ts_data                   (ftile_25gbe_rx_dma_ch1_rx_dma_fifo_0_in_ts_data),            //   input,   width = 96,                        .data
		.ftile_clk_clk                              (subsys_ftile_25gbe_1588_o_pll_clk_out_clk_clk),              //   input,    width = 1,               ftile_clk.clk
		.prefetcher_read_master_address             (rx_dma_ch1_prefetcher_read_master_address),                  //  output,   width = 37,  prefetcher_read_master.address
		.prefetcher_read_master_read                (rx_dma_ch1_prefetcher_read_master_read),                     //  output,    width = 1,                        .read
		.prefetcher_read_master_readdata            (rx_dma_ch1_prefetcher_read_master_readdata),                 //   input,  width = 128,                        .readdata
		.prefetcher_read_master_waitrequest         (rx_dma_ch1_prefetcher_read_master_waitrequest),              //   input,    width = 1,                        .waitrequest
		.prefetcher_read_master_readdatavalid       (rx_dma_ch1_prefetcher_read_master_readdatavalid),            //   input,    width = 1,                        .readdatavalid
		.prefetcher_read_master_burstcount          (rx_dma_ch1_prefetcher_read_master_burstcount),               //  output,    width = 3,                        .burstcount
		.prefetcher_write_master_address            (rx_dma_ch1_prefetcher_write_master_address),                 //  output,   width = 37, prefetcher_write_master.address
		.prefetcher_write_master_write              (rx_dma_ch1_prefetcher_write_master_write),                   //  output,    width = 1,                        .write
		.prefetcher_write_master_byteenable         (rx_dma_ch1_prefetcher_write_master_byteenable),              //  output,   width = 16,                        .byteenable
		.prefetcher_write_master_writedata          (rx_dma_ch1_prefetcher_write_master_writedata),               //  output,  width = 128,                        .writedata
		.prefetcher_write_master_waitrequest        (rx_dma_ch1_prefetcher_write_master_waitrequest),             //   input,    width = 1,                        .waitrequest
		.prefetcher_write_master_response           (rx_dma_ch1_prefetcher_write_master_response),                //   input,    width = 2,                        .response
		.prefetcher_write_master_writeresponsevalid (rx_dma_ch1_prefetcher_write_master_writeresponsevalid),      //   input,    width = 1,                        .writeresponsevalid
		.irq_irq                                    (rx_dma_ch1_irq_irq),                                         //  output,    width = 1,                     irq.irq
		.reset_reset_n                              (rx_dma_reset_bridge_out_reset_reset),                        //   input,    width = 1,                   reset.reset_n
		.write_master_address                       (rx_dma_ch1_write_master_address),                            //  output,   width = 37,            write_master.address
		.write_master_write                         (rx_dma_ch1_write_master_write),                              //  output,    width = 1,                        .write
		.write_master_byteenable                    (rx_dma_ch1_write_master_byteenable),                         //  output,   width = 16,                        .byteenable
		.write_master_writedata                     (rx_dma_ch1_write_master_writedata),                          //  output,  width = 128,                        .writedata
		.write_master_waitrequest                   (rx_dma_ch1_write_master_waitrequest),                        //   input,    width = 1,                        .waitrequest
		.write_master_burstcount                    (rx_dma_ch1_write_master_burstcount),                         //  output,    width = 5,                        .burstcount
		.write_master_response                      (rx_dma_ch1_write_master_response),                           //   input,    width = 2,                        .response
		.write_master_writeresponsevalid            (rx_dma_ch1_write_master_writeresponsevalid)                  //   input,    width = 1,                        .writeresponsevalid
	);

	subsys_ftile_25gbe_tx_dma #(
		.FP_WIDTH (FP_WIDTH)
	) ftile_25gbe_tx_dma_ch1 (
		.ts_chs_compl_0_clk_bus_in_clk              (ts_chs_compl_0_clk_bus_in_clk),                               //   input,    width = 1, ts_chs_compl_0_clk_bus_in.clk
		.ts_chs_compl_0_rst_bus_in_reset            (ts_chs_compl_0_rst_bus_in_reset),                             //   input,    width = 1, ts_chs_compl_0_rst_bus_in.reset
		.ts_chs_compl_0_i_ts_valid                  (ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_valid),            //   input,    width = 1,       ts_chs_compl_0_i_ts.valid
		.ts_chs_compl_0_i_ts_fingerprint            (ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_fingerprint),      //   input,   width = 20,                          .fingerprint
		.ts_chs_compl_0_i_ts_data                   (ftile_25gbe_tx_dma_ch1_ts_chs_compl_0_i_ts_data),             //   input,   width = 96,                          .data
		.dma_clk_clk                                (subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk),               //   input,    width = 1,                   dma_clk.clk
		.csr_waitrequest                            (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_waitrequest),    //  output,    width = 1,                       csr.waitrequest
		.csr_readdata                               (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_readdata),       //  output,   width = 32,                          .readdata
		.csr_readdatavalid                          (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_readdatavalid),  //  output,    width = 1,                          .readdatavalid
		.csr_burstcount                             (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_burstcount),     //   input,    width = 1,                          .burstcount
		.csr_writedata                              (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_writedata),      //   input,   width = 32,                          .writedata
		.csr_address                                (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_address),        //   input,    width = 6,                          .address
		.csr_write                                  (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_write),          //   input,    width = 1,                          .write
		.csr_read                                   (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_read),           //   input,    width = 1,                          .read
		.csr_byteenable                             (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_byteenable),     //   input,    width = 4,                          .byteenable
		.csr_debugaccess                            (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_debugaccess),    //   input,    width = 1,                          .debugaccess
		.tx_dma_fifo_0_out_st_ready                 (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_ready),           //   input,    width = 1,      tx_dma_fifo_0_out_st.ready
		.tx_dma_fifo_0_out_st_startofpacket         (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_startofpacket),   //  output,    width = 1,                          .startofpacket
		.tx_dma_fifo_0_out_st_valid                 (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_valid),           //  output,    width = 1,                          .valid
		.tx_dma_fifo_0_out_st_endofpacket           (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_endofpacket),     //  output,    width = 1,                          .endofpacket
		.tx_dma_fifo_0_out_st_data                  (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_data),            //  output,   width = 64,                          .data
		.tx_dma_fifo_0_out_st_empty                 (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_empty),           //  output,    width = 3,                          .empty
		.tx_dma_fifo_0_out_st_error                 (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_st_error),           //  output,    width = 1,                          .error
		.tx_dma_fifo_0_out_ts_req_valid             (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_valid),       //  output,    width = 1,  tx_dma_fifo_0_out_ts_req.valid
		.tx_dma_fifo_0_out_ts_req_fingerprint       (ftile_25gbe_tx_dma_ch1_tx_dma_fifo_0_out_ts_req_fingerprint), //  output,   width = 20,                          .fingerprint
		.ftile_clk_clk                              (subsys_ftile_25gbe_1588_o_pll_clk_out_clk_clk),               //   input,    width = 1,                 ftile_clk.clk
		.prefetcher_read_master_address             (tx_dma_ch1_prefetcher_read_master_address),                   //  output,   width = 37,    prefetcher_read_master.address
		.prefetcher_read_master_read                (tx_dma_ch1_prefetcher_read_master_read),                      //  output,    width = 1,                          .read
		.prefetcher_read_master_readdata            (tx_dma_ch1_prefetcher_read_master_readdata),                  //   input,  width = 128,                          .readdata
		.prefetcher_read_master_waitrequest         (tx_dma_ch1_prefetcher_read_master_waitrequest),               //   input,    width = 1,                          .waitrequest
		.prefetcher_read_master_readdatavalid       (tx_dma_ch1_prefetcher_read_master_readdatavalid),             //   input,    width = 1,                          .readdatavalid
		.prefetcher_read_master_burstcount          (tx_dma_ch1_prefetcher_read_master_burstcount),                //  output,    width = 3,                          .burstcount
		.prefetcher_write_master_address            (tx_dma_ch1_prefetcher_write_master_address),                  //  output,   width = 37,   prefetcher_write_master.address
		.prefetcher_write_master_write              (tx_dma_ch1_prefetcher_write_master_write),                    //  output,    width = 1,                          .write
		.prefetcher_write_master_byteenable         (tx_dma_ch1_prefetcher_write_master_byteenable),               //  output,   width = 16,                          .byteenable
		.prefetcher_write_master_writedata          (tx_dma_ch1_prefetcher_write_master_writedata),                //  output,  width = 128,                          .writedata
		.prefetcher_write_master_waitrequest        (tx_dma_ch1_prefetcher_write_master_waitrequest),              //   input,    width = 1,                          .waitrequest
		.prefetcher_write_master_response           (tx_dma_ch1_prefetcher_write_master_response),                 //   input,    width = 2,                          .response
		.prefetcher_write_master_writeresponsevalid (tx_dma_ch1_prefetcher_write_master_writeresponsevalid),       //   input,    width = 1,                          .writeresponsevalid
		.irq_irq                                    (tx_dma_ch1_irq_irq),                                          //  output,    width = 1,                       irq.irq
		.read_master_address                        (tx_dma_ch1_read_master_address),                              //  output,   width = 37,               read_master.address
		.read_master_read                           (tx_dma_ch1_read_master_read),                                 //  output,    width = 1,                          .read
		.read_master_byteenable                     (tx_dma_ch1_read_master_byteenable),                           //  output,   width = 16,                          .byteenable
		.read_master_readdata                       (tx_dma_ch1_read_master_readdata),                             //   input,  width = 128,                          .readdata
		.read_master_waitrequest                    (tx_dma_ch1_read_master_waitrequest),                          //   input,    width = 1,                          .waitrequest
		.read_master_readdatavalid                  (tx_dma_ch1_read_master_readdatavalid),                        //   input,    width = 1,                          .readdatavalid
		.read_master_burstcount                     (tx_dma_ch1_read_master_burstcount),                           //  output,    width = 5,                          .burstcount
		.reset_reset_n                              (~rst_controller_reset_out_reset)                              //   input,    width = 1,                     reset.reset_n
	);

	subsys_ftile_25gbe_1588_altera_mm_interconnect_1920_z5yfcuy mm_interconnect_0 (
		.subsys_ftile_25gbe_1588_csr_m0_address                                          (subsys_ftile_25gbe_1588_csr_m0_address),                     //   input,   width = 8,                                            subsys_ftile_25gbe_1588_csr_m0.address
		.subsys_ftile_25gbe_1588_csr_m0_waitrequest                                      (subsys_ftile_25gbe_1588_csr_m0_waitrequest),                 //  output,   width = 1,                                                                          .waitrequest
		.subsys_ftile_25gbe_1588_csr_m0_burstcount                                       (subsys_ftile_25gbe_1588_csr_m0_burstcount),                  //   input,   width = 1,                                                                          .burstcount
		.subsys_ftile_25gbe_1588_csr_m0_byteenable                                       (subsys_ftile_25gbe_1588_csr_m0_byteenable),                  //   input,   width = 4,                                                                          .byteenable
		.subsys_ftile_25gbe_1588_csr_m0_read                                             (subsys_ftile_25gbe_1588_csr_m0_read),                        //   input,   width = 1,                                                                          .read
		.subsys_ftile_25gbe_1588_csr_m0_readdata                                         (subsys_ftile_25gbe_1588_csr_m0_readdata),                    //  output,  width = 32,                                                                          .readdata
		.subsys_ftile_25gbe_1588_csr_m0_readdatavalid                                    (subsys_ftile_25gbe_1588_csr_m0_readdatavalid),               //  output,   width = 1,                                                                          .readdatavalid
		.subsys_ftile_25gbe_1588_csr_m0_write                                            (subsys_ftile_25gbe_1588_csr_m0_write),                       //   input,   width = 1,                                                                          .write
		.subsys_ftile_25gbe_1588_csr_m0_writedata                                        (subsys_ftile_25gbe_1588_csr_m0_writedata),                   //   input,  width = 32,                                                                          .writedata
		.subsys_ftile_25gbe_1588_csr_m0_debugaccess                                      (subsys_ftile_25gbe_1588_csr_m0_debugaccess),                 //   input,   width = 1,                                                                          .debugaccess
		.ftile_25gbe_tx_dma_ch1_csr_address                                              (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_address),       //  output,   width = 6,                                                ftile_25gbe_tx_dma_ch1_csr.address
		.ftile_25gbe_tx_dma_ch1_csr_write                                                (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_write),         //  output,   width = 1,                                                                          .write
		.ftile_25gbe_tx_dma_ch1_csr_read                                                 (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_read),          //  output,   width = 1,                                                                          .read
		.ftile_25gbe_tx_dma_ch1_csr_readdata                                             (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_readdata),      //   input,  width = 32,                                                                          .readdata
		.ftile_25gbe_tx_dma_ch1_csr_writedata                                            (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_writedata),     //  output,  width = 32,                                                                          .writedata
		.ftile_25gbe_tx_dma_ch1_csr_burstcount                                           (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_burstcount),    //  output,   width = 1,                                                                          .burstcount
		.ftile_25gbe_tx_dma_ch1_csr_byteenable                                           (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_byteenable),    //  output,   width = 4,                                                                          .byteenable
		.ftile_25gbe_tx_dma_ch1_csr_readdatavalid                                        (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_readdatavalid), //   input,   width = 1,                                                                          .readdatavalid
		.ftile_25gbe_tx_dma_ch1_csr_waitrequest                                          (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_waitrequest),   //   input,   width = 1,                                                                          .waitrequest
		.ftile_25gbe_tx_dma_ch1_csr_debugaccess                                          (mm_interconnect_0_ftile_25gbe_tx_dma_ch1_csr_debugaccess),   //  output,   width = 1,                                                                          .debugaccess
		.ftile_25gbe_rx_dma_ch1_csr_address                                              (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_address),       //  output,   width = 6,                                                ftile_25gbe_rx_dma_ch1_csr.address
		.ftile_25gbe_rx_dma_ch1_csr_write                                                (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_write),         //  output,   width = 1,                                                                          .write
		.ftile_25gbe_rx_dma_ch1_csr_read                                                 (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_read),          //  output,   width = 1,                                                                          .read
		.ftile_25gbe_rx_dma_ch1_csr_readdata                                             (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_readdata),      //   input,  width = 32,                                                                          .readdata
		.ftile_25gbe_rx_dma_ch1_csr_writedata                                            (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_writedata),     //  output,  width = 32,                                                                          .writedata
		.ftile_25gbe_rx_dma_ch1_csr_burstcount                                           (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_burstcount),    //  output,   width = 1,                                                                          .burstcount
		.ftile_25gbe_rx_dma_ch1_csr_byteenable                                           (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_byteenable),    //  output,   width = 4,                                                                          .byteenable
		.ftile_25gbe_rx_dma_ch1_csr_readdatavalid                                        (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_readdatavalid), //   input,   width = 1,                                                                          .readdatavalid
		.ftile_25gbe_rx_dma_ch1_csr_waitrequest                                          (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_waitrequest),   //   input,   width = 1,                                                                          .waitrequest
		.ftile_25gbe_rx_dma_ch1_csr_debugaccess                                          (mm_interconnect_0_ftile_25gbe_rx_dma_ch1_csr_debugaccess),   //  output,   width = 1,                                                                          .debugaccess
		.subsys_ftile_25gbe_1588_csr_reset_reset_bridge_in_reset_reset                   (~subsys_ftile_25gbe_1588_reset_out_reset_reset),             //   input,   width = 1,                   subsys_ftile_25gbe_1588_csr_reset_reset_bridge_in_reset.reset
		.ftile_25gbe_tx_dma_ch1_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                             //   input,   width = 1,                        ftile_25gbe_tx_dma_ch1_reset_reset_bridge_in_reset.reset
		.ftile_25gbe_rx_dma_ch1_reset_reset_bridge_in_reset_reset                        (~rx_dma_reset_bridge_out_reset_reset),                       //   input,   width = 1,                        ftile_25gbe_rx_dma_ch1_reset_reset_bridge_in_reset.reset
		.subsys_ftile_25gbe_1588_csr_m0_translator_reset_reset_bridge_in_reset_reset     (~subsys_ftile_25gbe_1588_reset_out_reset_reset),             //   input,   width = 1,     subsys_ftile_25gbe_1588_csr_m0_translator_reset_reset_bridge_in_reset.reset
		.ftile_25gbe_tx_dma_ch1_csr_agent_rsp_fifo_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             //   input,   width = 1, ftile_25gbe_tx_dma_ch1_csr_agent_rsp_fifo_clk_reset_reset_bridge_in_reset.reset
		.ftile_25gbe_rx_dma_ch1_csr_agent_rsp_fifo_clk_reset_reset_bridge_in_reset_reset (~rx_dma_reset_bridge_out_reset_reset),                       //   input,   width = 1, ftile_25gbe_rx_dma_ch1_csr_agent_rsp_fifo_clk_reset_reset_bridge_in_reset.reset
		.subsys_ftile_25gbe_1588_csrclk_out_clk_clk                                      (subsys_ftile_25gbe_1588_csrclk_out_clk_clk),                 //   input,   width = 1,                                    subsys_ftile_25gbe_1588_csrclk_out_clk.clk
		.subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk                                   (subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk)               //   input,   width = 1,                                 subsys_ftile_25gbe_1588_dmaclkout_out_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~subsys_ftile_25gbe_1588_reset_out_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (subsys_ftile_25gbe_1588_dmaclkout_out_clk_clk),  //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                 //  output,  width = 1, reset_out.reset
		.reset_req      (),                                               // (terminated),                       
		.reset_req_in0  (1'b0),                                           // (terminated),                       
		.reset_in1      (1'b0),                                           // (terminated),                       
		.reset_req_in1  (1'b0),                                           // (terminated),                       
		.reset_in2      (1'b0),                                           // (terminated),                       
		.reset_req_in2  (1'b0),                                           // (terminated),                       
		.reset_in3      (1'b0),                                           // (terminated),                       
		.reset_req_in3  (1'b0),                                           // (terminated),                       
		.reset_in4      (1'b0),                                           // (terminated),                       
		.reset_req_in4  (1'b0),                                           // (terminated),                       
		.reset_in5      (1'b0),                                           // (terminated),                       
		.reset_req_in5  (1'b0),                                           // (terminated),                       
		.reset_in6      (1'b0),                                           // (terminated),                       
		.reset_req_in6  (1'b0),                                           // (terminated),                       
		.reset_in7      (1'b0),                                           // (terminated),                       
		.reset_req_in7  (1'b0),                                           // (terminated),                       
		.reset_in8      (1'b0),                                           // (terminated),                       
		.reset_req_in8  (1'b0),                                           // (terminated),                       
		.reset_in9      (1'b0),                                           // (terminated),                       
		.reset_req_in9  (1'b0),                                           // (terminated),                       
		.reset_in10     (1'b0),                                           // (terminated),                       
		.reset_req_in10 (1'b0),                                           // (terminated),                       
		.reset_in11     (1'b0),                                           // (terminated),                       
		.reset_req_in11 (1'b0),                                           // (terminated),                       
		.reset_in12     (1'b0),                                           // (terminated),                       
		.reset_req_in12 (1'b0),                                           // (terminated),                       
		.reset_in13     (1'b0),                                           // (terminated),                       
		.reset_req_in13 (1'b0),                                           // (terminated),                       
		.reset_in14     (1'b0),                                           // (terminated),                       
		.reset_req_in14 (1'b0),                                           // (terminated),                       
		.reset_in15     (1'b0),                                           // (terminated),                       
		.reset_req_in15 (1'b0)                                            // (terminated),                       
	);

endmodule
